module Test( // @[when_test.py:15:when_test.fir@2.2]
  input         clock, // @[rawmodule.py:100:when_test.fir@3.4]
  input         reset, // @[rawmodule.py:101:when_test.fir@4.4]
  input  [31:0] io_a, // @[when_test.py:6:when_test.fir@5.4]
  input  [31:0] io_b, // @[when_test.py:6:when_test.fir@5.4]
  input  [3:0]  io_sig, // @[when_test.py:6:when_test.fir@5.4]
  output [31:0] io_out // @[when_test.py:6:when_test.fir@5.4]
);
  wire  _T_9; // @[when_test.py:18:when_test.fir@8.4]
  wire  _T_12; // @[when_test.py:20:when_test.fir@13.6]
  wire  _T_13; // @[when_test.py:20:when_test.fir@14.6]
  wire  _T_14; // @[when_test.py:20:when_test.fir@15.6]
  wire  _T_17; // @[when_test.py:22:when_test.fir@20.8]
  wire  _T_18; // @[when_test.py:22:when_test.fir@21.8]
  wire  _T_19; // @[when_test.py:22:when_test.fir@22.8]
  wire [63:0] _T_20; // @[when_test.py:23:when_test.fir@24.10]
  wire [3:0] _T_21; // @[when_test.py:24:when_test.fir@28.10]
  wire  _T_23; // @[when_test.py:24:when_test.fir@30.10]
  wire [31:0] _T_24; // @[when_test.py:25:when_test.fir@32.12]
  wire  _T_25; // @[when_test.py:26:when_test.fir@36.12]
  wire  _T_26; // @[when_test.py:26:when_test.fir@37.12]
  wire  _T_27; // @[when_test.py:26:when_test.fir@38.12]
  wire [31:0] _T_28; // @[when_test.py:27:when_test.fir@40.14]
  wire [31:0] _T_29; // @[when_test.py:29:when_test.fir@44.14]
  wire [31:0] _GEN_0; // @[when_test.py:26:when_test.fir@39.12]
  wire [31:0] _GEN_1; // @[when_test.py:24:when_test.fir@31.10]
  wire [63:0] _GEN_2; // @[when_test.py:22:when_test.fir@23.8]
  wire  _T_30; // @[when_test.py:30:when_test.fir@51.8]
  wire  _T_31; // @[when_test.py:30:when_test.fir@52.8]
  wire  _T_32; // @[when_test.py:30:when_test.fir@53.8]
  wire [31:0] _T_33; // @[when_test.py:31:when_test.fir@55.10]
  wire  _T_34; // @[when_test.py:32:when_test.fir@59.10]
  wire  _T_35; // @[when_test.py:32:when_test.fir@60.10]
  wire  _T_36; // @[when_test.py:32:when_test.fir@61.10]
  wire [31:0] _GEN_9; // @[when_test.py:33:when_test.fir@63.12]
  wire [31:0] _T_37; // @[when_test.py:33:when_test.fir@63.12]
  wire  _T_38; // @[when_test.py:35:when_test.fir@67.12]
  wire [31:0] _GEN_3; // @[when_test.py:32:when_test.fir@62.10]
  wire [31:0] _GEN_4; // @[when_test.py:30:when_test.fir@54.8]
  wire [63:0] _GEN_5; // @[when_test.py:20:when_test.fir@16.6]
  wire  _T_39; // @[when_test.py:36:when_test.fir@74.6]
  wire  _T_40; // @[when_test.py:36:when_test.fir@75.6]
  wire  _T_41; // @[when_test.py:36:when_test.fir@76.6]
  wire  _T_42; // @[when_test.py:37:when_test.fir@78.8]
  wire  _T_43; // @[when_test.py:38:when_test.fir@82.8]
  wire  _T_44; // @[when_test.py:38:when_test.fir@83.8]
  wire  _T_45; // @[when_test.py:38:when_test.fir@84.8]
  wire  _T_46; // @[when_test.py:39:when_test.fir@86.10]
  wire  _T_47; // @[when_test.py:41:when_test.fir@90.10]
  wire  _GEN_6; // @[when_test.py:38:when_test.fir@85.8]
  wire  _GEN_7; // @[when_test.py:36:when_test.fir@77.6]
  wire [63:0] _GEN_8; // @[when_test.py:18:when_test.fir@10.4]
  assign _T_9 = io_sig < 4'h1; // @[when_test.py:18:when_test.fir@8.4]
  assign _T_12 = io_sig >= 4'h1; // @[when_test.py:20:when_test.fir@13.6]
  assign _T_13 = io_sig < 4'h2; // @[when_test.py:20:when_test.fir@14.6]
  assign _T_14 = _T_12 & _T_13; // @[when_test.py:20:when_test.fir@15.6]
  assign _T_17 = io_sig >= 4'h2; // @[when_test.py:22:when_test.fir@20.8]
  assign _T_18 = io_sig < 4'h3; // @[when_test.py:22:when_test.fir@21.8]
  assign _T_19 = _T_17 & _T_18; // @[when_test.py:22:when_test.fir@22.8]
  assign _T_20 = io_a * io_b; // @[when_test.py:23:when_test.fir@24.10]
  assign _T_21 = 4'h3 & io_sig; // @[when_test.py:24:when_test.fir@28.10]
  assign _T_23 = _T_21 < 4'h4; // @[when_test.py:24:when_test.fir@30.10]
  assign _T_24 = io_a / io_b; // @[when_test.py:25:when_test.fir@32.12]
  assign _T_25 = io_sig >= 4'h4; // @[when_test.py:26:when_test.fir@36.12]
  assign _T_26 = io_sig < 4'h5; // @[when_test.py:26:when_test.fir@37.12]
  assign _T_27 = _T_25 & _T_26; // @[when_test.py:26:when_test.fir@38.12]
  assign _T_28 = io_a & io_b; // @[when_test.py:27:when_test.fir@40.14]
  assign _T_29 = io_a | io_b; // @[when_test.py:29:when_test.fir@44.14]
  assign _GEN_0 = _T_27 ? _T_28 : _T_29; // @[when_test.py:26:when_test.fir@39.12]
  assign _GEN_1 = _T_23 ? _T_24 : _GEN_0; // @[when_test.py:24:when_test.fir@31.10]
  assign _GEN_2 = _T_19 ? _T_20 : {{32'd0}, _GEN_1}; // @[when_test.py:22:when_test.fir@23.8]
  assign _T_30 = io_sig >= 4'h5; // @[when_test.py:30:when_test.fir@51.8]
  assign _T_31 = io_sig < 4'h6; // @[when_test.py:30:when_test.fir@52.8]
  assign _T_32 = _T_30 & _T_31; // @[when_test.py:30:when_test.fir@53.8]
  assign _T_33 = io_a ^ io_b; // @[when_test.py:31:when_test.fir@55.10]
  assign _T_34 = io_sig >= 4'h6; // @[when_test.py:32:when_test.fir@59.10]
  assign _T_35 = io_sig < 4'h7; // @[when_test.py:32:when_test.fir@60.10]
  assign _T_36 = _T_34 & _T_35; // @[when_test.py:32:when_test.fir@61.10]
  assign _GEN_9 = io_a % io_b; // @[when_test.py:33:when_test.fir@63.12]
  assign _T_37 = _GEN_9[31:0]; // @[when_test.py:33:when_test.fir@63.12]
  assign _T_38 = io_a == io_b; // @[when_test.py:35:when_test.fir@67.12]
  assign _GEN_3 = _T_36 ? _T_37 : {{31'd0}, _T_38}; // @[when_test.py:32:when_test.fir@62.10]
  assign _GEN_4 = _T_32 ? _T_33 : _GEN_3; // @[when_test.py:30:when_test.fir@54.8]
  assign _GEN_5 = _T_14 ? _GEN_2 : {{32'd0}, _GEN_4}; // @[when_test.py:20:when_test.fir@16.6]
  assign _T_39 = io_sig >= 4'h7; // @[when_test.py:36:when_test.fir@74.6]
  assign _T_40 = io_sig < 4'h8; // @[when_test.py:36:when_test.fir@75.6]
  assign _T_41 = _T_39 & _T_40; // @[when_test.py:36:when_test.fir@76.6]
  assign _T_42 = io_a != io_b; // @[when_test.py:37:when_test.fir@78.8]
  assign _T_43 = io_sig >= 4'h8; // @[when_test.py:38:when_test.fir@82.8]
  assign _T_44 = io_sig < 4'h9; // @[when_test.py:38:when_test.fir@83.8]
  assign _T_45 = _T_43 & _T_44; // @[when_test.py:38:when_test.fir@84.8]
  assign _T_46 = io_a < io_b; // @[when_test.py:39:when_test.fir@86.10]
  assign _T_47 = io_a > io_b; // @[when_test.py:41:when_test.fir@90.10]
  assign _GEN_6 = _T_45 ? _T_46 : _T_47; // @[when_test.py:38:when_test.fir@85.8]
  assign _GEN_7 = _T_41 ? _T_42 : _GEN_6; // @[when_test.py:36:when_test.fir@77.6]
  assign _GEN_8 = _T_9 ? _GEN_5 : {{63'd0}, _GEN_7}; // @[when_test.py:18:when_test.fir@10.4]
  assign io_out = _GEN_8[31:0]; // @[when_test.py:19:when_test.fir@12.6 when_test.py:21:when_test.fir@19.8 when_test.py:23:when_test.fir@25.10 when_test.py:25:when_test.fir@33.12 when_test.py:27:when_test.fir@41.14 when_test.py:29:when_test.fir@45.14 when_test.py:31:when_test.fir@56.10 when_test.py:33:when_test.fir@64.12 when_test.py:35:when_test.fir@68.12 when_test.py:37:when_test.fir@79.8 when_test.py:39:when_test.fir@87.10 when_test.py:41:when_test.fir@91.10]
endmodule
