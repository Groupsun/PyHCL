module Datapath( // @[datapath.py:94:datapath.fir@2.2]
  input         clock, // @[rawmodule.py:100:datapath.fir@3.4]
  input         reset, // @[rawmodule.py:101:datapath.fir@4.4]
  input  [31:0] io_if_io_if_pc, // @[datapath.py:84:datapath.fir@5.4]
  input  [1:0]  io_if_io_PC_Sel, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_if_io_new_addr, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_if_io_pc_recover, // @[datapath.py:84:datapath.fir@5.4]
  output [31:0] io_if_io_if_new_pc, // @[datapath.py:84:datapath.fir@5.4]
  output [31:0] io_if_io_if_pc_4, // @[datapath.py:84:datapath.fir@5.4]
  input         io_id_io_Bubble, // @[datapath.py:84:datapath.fir@5.4]
  input         io_id_io_ctrl_in_Reg_Write, // @[datapath.py:84:datapath.fir@5.4]
  input  [2:0]  io_id_io_ctrl_in_Imm_Sel, // @[datapath.py:84:datapath.fir@5.4]
  input         io_id_io_ctrl_in_ALU_Src, // @[datapath.py:84:datapath.fir@5.4]
  input  [4:0]  io_id_io_ctrl_in_ALUOp, // @[datapath.py:84:datapath.fir@5.4]
  input         io_id_io_ctrl_in_Branch, // @[datapath.py:84:datapath.fir@5.4]
  input         io_id_io_ctrl_in_Branch_Src, // @[datapath.py:84:datapath.fir@5.4]
  input         io_id_io_ctrl_in_Mem_Read, // @[datapath.py:84:datapath.fir@5.4]
  input         io_id_io_ctrl_in_Mem_Write, // @[datapath.py:84:datapath.fir@5.4]
  input  [1:0]  io_id_io_ctrl_in_Data_Size, // @[datapath.py:84:datapath.fir@5.4]
  input         io_id_io_ctrl_in_Load_Type, // @[datapath.py:84:datapath.fir@5.4]
  input  [2:0]  io_id_io_ctrl_in_Mem_to_Reg, // @[datapath.py:84:datapath.fir@5.4]
  input         io_id_io_ctrl_in_Jump_Type, // @[datapath.py:84:datapath.fir@5.4]
  output        io_id_io_ctrl_out_Reg_Write, // @[datapath.py:84:datapath.fir@5.4]
  output [2:0]  io_id_io_ctrl_out_Imm_Sel, // @[datapath.py:84:datapath.fir@5.4]
  output        io_id_io_ctrl_out_ALU_Src, // @[datapath.py:84:datapath.fir@5.4]
  output [4:0]  io_id_io_ctrl_out_ALUOp, // @[datapath.py:84:datapath.fir@5.4]
  output        io_id_io_ctrl_out_Branch, // @[datapath.py:84:datapath.fir@5.4]
  output        io_id_io_ctrl_out_Branch_Src, // @[datapath.py:84:datapath.fir@5.4]
  output        io_id_io_ctrl_out_Mem_Read, // @[datapath.py:84:datapath.fir@5.4]
  output        io_id_io_ctrl_out_Mem_Write, // @[datapath.py:84:datapath.fir@5.4]
  output [1:0]  io_id_io_ctrl_out_Data_Size, // @[datapath.py:84:datapath.fir@5.4]
  output        io_id_io_ctrl_out_Load_Type, // @[datapath.py:84:datapath.fir@5.4]
  output [2:0]  io_id_io_ctrl_out_Mem_to_Reg, // @[datapath.py:84:datapath.fir@5.4]
  output        io_id_io_ctrl_out_Jump_Type, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_ex_io_ex_rs1_out, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_ex_io_ex_rs2_out, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_ex_io_ex_imm, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_ex_io_ex_pc, // @[datapath.py:84:datapath.fir@5.4]
  input         io_ex_io_ex_ALU_Src, // @[datapath.py:84:datapath.fir@5.4]
  input         io_ex_io_ex_Branch, // @[datapath.py:84:datapath.fir@5.4]
  input         io_ex_io_ex_alu_conflag, // @[datapath.py:84:datapath.fir@5.4]
  input         io_ex_io_ex_Branch_Src, // @[datapath.py:84:datapath.fir@5.4]
  input         io_ex_io_ex_Jump_Type, // @[datapath.py:84:datapath.fir@5.4]
  input  [2:0]  io_ex_io_ex_Imm_Sel, // @[datapath.py:84:datapath.fir@5.4]
  input  [1:0]  io_ex_io_Forward_A, // @[datapath.py:84:datapath.fir@5.4]
  input  [1:0]  io_ex_io_Forward_B, // @[datapath.py:84:datapath.fir@5.4]
  output [31:0] io_ex_io_alu_a_src, // @[datapath.py:84:datapath.fir@5.4]
  output [31:0] io_ex_io_alu_b_src, // @[datapath.py:84:datapath.fir@5.4]
  output [31:0] io_ex_io_ex_aui_pc, // @[datapath.py:84:datapath.fir@5.4]
  output [31:0] io_ex_io_forward_rs2_out, // @[datapath.py:84:datapath.fir@5.4]
  output        io_ex_io_PC_Src, // @[datapath.py:84:datapath.fir@5.4]
  output [31:0] io_ex_io_branch_addr, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_mem_io_mem_rs2_out, // @[datapath.py:84:datapath.fir@5.4]
  input         io_mem_io_MemWrite_Src, // @[datapath.py:84:datapath.fir@5.4]
  input  [2:0]  io_mem_io_mem_Mem_to_Reg, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_mem_io_mem_alu_sum, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_mem_io_mem_pc_4, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_mem_io_mem_imm, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_mem_io_mem_aui_pc, // @[datapath.py:84:datapath.fir@5.4]
  output [31:0] io_mem_io_mem_writedata, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_wb_io_wb_alu_sum, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_wb_io_wb_dataout, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_wb_io_wb_pc_4, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_wb_io_wb_imm, // @[datapath.py:84:datapath.fir@5.4]
  input  [31:0] io_wb_io_wb_aui_pc, // @[datapath.py:84:datapath.fir@5.4]
  input  [2:0]  io_wb_io_wb_Mem_to_Reg, // @[datapath.py:84:datapath.fir@5.4]
  output [31:0] io_wb_io_wb_reg_writedata // @[datapath.py:84:datapath.fir@5.4]
);
  wire  _T_82; // @[datapath.py:103:datapath.fir@7.4]
  wire  _T_84; // @[datapath.py:103:datapath.fir@9.4]
  wire [32:0] _T_85; // @[datapath.py:105:datapath.fir@10.4]
  wire [32:0] _T_86; // @[datapath.py:108:datapath.fir@12.4]
  wire [32:0] _T_87; // @[datapath.py:108:datapath.fir@13.4]
  wire [31:0] _T_89; // @[datapath.py:109:datapath.fir@15.4]
  wire [32:0] _T_90; // @[datapath.py:110:datapath.fir@16.4]
  wire [32:0] _GEN_0; // @[datapath.py:110:datapath.fir@17.4]
  wire [33:0] _T_91; // @[datapath.py:110:datapath.fir@17.4]
  wire [32:0] _T_94; // @[datapath.py:112:datapath.fir@20.4]
  wire  _T_96; // @[datapath.py:116:datapath.fir@24.4]
  wire  _T_100; // @[mux.py:72:datapath.fir@29.4]
  wire [31:0] _T_101; // @[datapath.py:123:datapath.fir@30.4]
  wire  _T_102; // @[mux.py:72:datapath.fir@31.4]
  wire [31:0] _T_103; // @[datapath.py:123:datapath.fir@32.4]
  wire  _T_104; // @[mux.py:72:datapath.fir@33.4]
  wire [32:0] _T_105; // @[datapath.py:123:datapath.fir@34.4]
  wire  _T_130; // @[mux.py:72:datapath.fir@72.4]
  wire [31:0] _T_131; // @[datapath.py:146:datapath.fir@73.4]
  wire  _T_132; // @[mux.py:72:datapath.fir@74.4]
  wire [31:0] _T_133; // @[datapath.py:146:datapath.fir@75.4]
  wire  _T_134; // @[mux.py:72:datapath.fir@76.4]
  wire [31:0] _T_135; // @[datapath.py:146:datapath.fir@77.4]
  wire  _T_136; // @[mux.py:72:datapath.fir@78.4]
  wire [31:0] _T_137; // @[datapath.py:146:datapath.fir@79.4]
  wire  _T_138; // @[mux.py:72:datapath.fir@80.4]
  wire [31:0] _T_139; // @[datapath.py:152:datapath.fir@81.4]
  wire  _T_140; // @[mux.py:72:datapath.fir@82.4]
  wire [31:0] _T_141; // @[datapath.py:152:datapath.fir@83.4]
  wire  _T_142; // @[mux.py:72:datapath.fir@84.4]
  wire  _T_144; // @[mux.py:72:datapath.fir@87.4]
  wire [31:0] _T_145; // @[datapath.py:158:datapath.fir@88.4]
  wire  _T_146; // @[mux.py:72:datapath.fir@89.4]
  wire [31:0] _T_147; // @[datapath.py:158:datapath.fir@90.4]
  wire  _T_148; // @[mux.py:72:datapath.fir@91.4]
  wire [31:0] _T_149; // @[datapath.py:158:datapath.fir@92.4]
  wire  _T_154; // @[mux.py:72:datapath.fir@100.4]
  wire [31:0] _T_155; // @[datapath.py:180:datapath.fir@101.4]
  wire  _T_156; // @[mux.py:72:datapath.fir@102.4]
  wire [31:0] _T_157; // @[datapath.py:180:datapath.fir@103.4]
  wire  _T_158; // @[mux.py:72:datapath.fir@104.4]
  wire [31:0] _T_159; // @[datapath.py:180:datapath.fir@105.4]
  wire  _T_160; // @[mux.py:72:datapath.fir@106.4]
  wire [31:0] _T_161; // @[datapath.py:180:datapath.fir@107.4]
  wire  _T_162; // @[mux.py:72:datapath.fir@108.4]
  assign _T_82 = io_ex_io_ex_Imm_Sel == 3'h2; // @[datapath.py:103:datapath.fir@7.4]
  assign _T_84 = _T_82 & io_ex_io_ex_Jump_Type; // @[datapath.py:103:datapath.fir@9.4]
  assign _T_85 = io_if_io_if_pc + 32'h4; // @[datapath.py:105:datapath.fir@10.4]
  assign _T_86 = {io_ex_io_ex_imm, 1'h0}; // @[datapath.py:108:datapath.fir@12.4]
  assign _T_87 = _T_84 ? {{1'd0}, io_ex_io_ex_imm} : _T_86; // @[datapath.py:108:datapath.fir@13.4]
  assign _T_89 = io_ex_io_ex_Branch_Src ? io_ex_io_alu_a_src : io_ex_io_ex_pc; // @[datapath.py:109:datapath.fir@15.4]
  assign _T_90 = $unsigned(_T_87); // @[datapath.py:110:datapath.fir@16.4]
  assign _GEN_0 = {{1'd0}, _T_89}; // @[datapath.py:110:datapath.fir@17.4]
  assign _T_91 = _GEN_0 + _T_90; // @[datapath.py:110:datapath.fir@17.4]
  assign _T_94 = _T_89 + io_ex_io_ex_imm; // @[datapath.py:112:datapath.fir@20.4]
  assign _T_96 = io_ex_io_ex_Jump_Type ? 1'h1 : io_ex_io_ex_alu_conflag; // @[datapath.py:116:datapath.fir@24.4]
  assign _T_100 = io_if_io_PC_Sel == 2'h1; // @[mux.py:72:datapath.fir@29.4]
  assign _T_101 = _T_100 ? io_if_io_pc_recover : 32'h0; // @[datapath.py:123:datapath.fir@30.4]
  assign _T_102 = io_if_io_PC_Sel == 2'h2; // @[mux.py:72:datapath.fir@31.4]
  assign _T_103 = _T_102 ? io_if_io_new_addr : _T_101; // @[datapath.py:123:datapath.fir@32.4]
  assign _T_104 = io_if_io_PC_Sel == 2'h0; // @[mux.py:72:datapath.fir@33.4]
  assign _T_105 = _T_104 ? _T_85 : {{1'd0}, _T_103}; // @[datapath.py:123:datapath.fir@34.4]
  assign _T_130 = io_mem_io_mem_Mem_to_Reg == 3'h4; // @[mux.py:72:datapath.fir@72.4]
  assign _T_131 = _T_130 ? io_mem_io_mem_aui_pc : 32'h0; // @[datapath.py:146:datapath.fir@73.4]
  assign _T_132 = io_mem_io_mem_Mem_to_Reg == 3'h3; // @[mux.py:72:datapath.fir@74.4]
  assign _T_133 = _T_132 ? io_mem_io_mem_imm : _T_131; // @[datapath.py:146:datapath.fir@75.4]
  assign _T_134 = io_mem_io_mem_Mem_to_Reg == 3'h2; // @[mux.py:72:datapath.fir@76.4]
  assign _T_135 = _T_134 ? io_mem_io_mem_pc_4 : _T_133; // @[datapath.py:146:datapath.fir@77.4]
  assign _T_136 = io_mem_io_mem_Mem_to_Reg == 3'h0; // @[mux.py:72:datapath.fir@78.4]
  assign _T_137 = _T_136 ? io_mem_io_mem_alu_sum : _T_135; // @[datapath.py:146:datapath.fir@79.4]
  assign _T_138 = io_ex_io_Forward_A == 2'h2; // @[mux.py:72:datapath.fir@80.4]
  assign _T_139 = _T_138 ? _T_137 : io_ex_io_ex_rs1_out; // @[datapath.py:152:datapath.fir@81.4]
  assign _T_140 = io_ex_io_Forward_A == 2'h1; // @[mux.py:72:datapath.fir@82.4]
  assign _T_141 = _T_140 ? io_wb_io_wb_reg_writedata : _T_139; // @[datapath.py:152:datapath.fir@83.4]
  assign _T_142 = io_ex_io_Forward_A == 2'h0; // @[mux.py:72:datapath.fir@84.4]
  assign _T_144 = io_ex_io_Forward_B == 2'h2; // @[mux.py:72:datapath.fir@87.4]
  assign _T_145 = _T_144 ? _T_137 : io_ex_io_ex_rs2_out; // @[datapath.py:158:datapath.fir@88.4]
  assign _T_146 = io_ex_io_Forward_B == 2'h1; // @[mux.py:72:datapath.fir@89.4]
  assign _T_147 = _T_146 ? io_wb_io_wb_reg_writedata : _T_145; // @[datapath.py:158:datapath.fir@90.4]
  assign _T_148 = io_ex_io_Forward_B == 2'h0; // @[mux.py:72:datapath.fir@91.4]
  assign _T_149 = _T_148 ? io_ex_io_ex_rs2_out : _T_147; // @[datapath.py:158:datapath.fir@92.4]
  assign _T_154 = io_wb_io_wb_Mem_to_Reg == 3'h4; // @[mux.py:72:datapath.fir@100.4]
  assign _T_155 = _T_154 ? io_wb_io_wb_aui_pc : io_wb_io_wb_alu_sum; // @[datapath.py:180:datapath.fir@101.4]
  assign _T_156 = io_wb_io_wb_Mem_to_Reg == 3'h3; // @[mux.py:72:datapath.fir@102.4]
  assign _T_157 = _T_156 ? io_wb_io_wb_imm : _T_155; // @[datapath.py:180:datapath.fir@103.4]
  assign _T_158 = io_wb_io_wb_Mem_to_Reg == 3'h2; // @[mux.py:72:datapath.fir@104.4]
  assign _T_159 = _T_158 ? io_wb_io_wb_pc_4 : _T_157; // @[datapath.py:180:datapath.fir@105.4]
  assign _T_160 = io_wb_io_wb_Mem_to_Reg == 3'h1; // @[mux.py:72:datapath.fir@106.4]
  assign _T_161 = _T_160 ? io_wb_io_wb_dataout : _T_159; // @[datapath.py:180:datapath.fir@107.4]
  assign _T_162 = io_wb_io_wb_Mem_to_Reg == 3'h0; // @[mux.py:72:datapath.fir@108.4]
  assign io_if_io_if_new_pc = _T_105[31:0]; // @[datapath.py:123:datapath.fir@35.4]
  assign io_if_io_if_pc_4 = _T_85[31:0]; // @[datapath.py:106:datapath.fir@11.4]
  assign io_id_io_ctrl_out_Reg_Write = io_id_io_Bubble ? 1'h0 : io_id_io_ctrl_in_Reg_Write; // @[datapath.py:135:datapath.fir@38.4]
  assign io_id_io_ctrl_out_Imm_Sel = io_id_io_Bubble ? 3'h0 : io_id_io_ctrl_in_Imm_Sel; // @[datapath.py:135:datapath.fir@41.4]
  assign io_id_io_ctrl_out_ALU_Src = io_id_io_Bubble ? 1'h0 : io_id_io_ctrl_in_ALU_Src; // @[datapath.py:135:datapath.fir@44.4]
  assign io_id_io_ctrl_out_ALUOp = io_id_io_Bubble ? 5'h0 : io_id_io_ctrl_in_ALUOp; // @[datapath.py:135:datapath.fir@47.4]
  assign io_id_io_ctrl_out_Branch = io_id_io_Bubble ? 1'h0 : io_id_io_ctrl_in_Branch; // @[datapath.py:135:datapath.fir@50.4]
  assign io_id_io_ctrl_out_Branch_Src = io_id_io_Bubble ? 1'h0 : io_id_io_ctrl_in_Branch_Src; // @[datapath.py:135:datapath.fir@53.4]
  assign io_id_io_ctrl_out_Mem_Read = io_id_io_Bubble ? 1'h0 : io_id_io_ctrl_in_Mem_Read; // @[datapath.py:135:datapath.fir@56.4]
  assign io_id_io_ctrl_out_Mem_Write = io_id_io_Bubble ? 1'h0 : io_id_io_ctrl_in_Mem_Write; // @[datapath.py:135:datapath.fir@59.4]
  assign io_id_io_ctrl_out_Data_Size = io_id_io_Bubble ? 2'h0 : io_id_io_ctrl_in_Data_Size; // @[datapath.py:135:datapath.fir@62.4]
  assign io_id_io_ctrl_out_Load_Type = io_id_io_Bubble ? 1'h0 : io_id_io_ctrl_in_Load_Type; // @[datapath.py:135:datapath.fir@65.4]
  assign io_id_io_ctrl_out_Mem_to_Reg = io_id_io_Bubble ? 3'h0 : io_id_io_ctrl_in_Mem_to_Reg; // @[datapath.py:135:datapath.fir@68.4]
  assign io_id_io_ctrl_out_Jump_Type = io_id_io_Bubble ? 1'h0 : io_id_io_ctrl_in_Jump_Type; // @[datapath.py:135:datapath.fir@71.4]
  assign io_ex_io_alu_a_src = _T_142 ? io_ex_io_ex_rs1_out : _T_141; // @[datapath.py:152:datapath.fir@86.4]
  assign io_ex_io_alu_b_src = io_ex_io_ex_ALU_Src ? io_ex_io_ex_imm : _T_149; // @[datapath.py:162:datapath.fir@95.4]
  assign io_ex_io_ex_aui_pc = _T_94[31:0]; // @[datapath.py:112:datapath.fir@21.4]
  assign io_ex_io_forward_rs2_out = _T_148 ? io_ex_io_ex_rs2_out : _T_147; // @[datapath.py:163:datapath.fir@96.4]
  assign io_ex_io_PC_Src = _T_96 & io_ex_io_ex_Branch; // @[datapath.py:118:datapath.fir@28.4]
  assign io_ex_io_branch_addr = _T_91[31:0]; // @[datapath.py:113:datapath.fir@22.4]
  assign io_mem_io_mem_writedata = io_mem_io_MemWrite_Src ? io_wb_io_wb_reg_writedata : io_mem_io_mem_rs2_out; // @[datapath.py:169:datapath.fir@99.4]
  assign io_wb_io_wb_reg_writedata = _T_162 ? io_wb_io_wb_alu_sum : _T_161; // @[datapath.py:180:datapath.fir@110.4]
endmodule
