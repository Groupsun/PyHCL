module Control( // @[control.py:92:Control.fir@2.2]
  input         clock, // @[rawmodule.py:100:Control.fir@3.4]
  input         reset, // @[rawmodule.py:101:Control.fir@4.4]
  input  [31:0] io_inst, // @[control.py:85:Control.fir@5.4]
  output        io_ctrl_Reg_Write, // @[control.py:85:Control.fir@5.4]
  output [2:0]  io_ctrl_Imm_Sel, // @[control.py:85:Control.fir@5.4]
  output        io_ctrl_ALU_Src, // @[control.py:85:Control.fir@5.4]
  output [4:0]  io_ctrl_ALUOp, // @[control.py:85:Control.fir@5.4]
  output        io_ctrl_Branch, // @[control.py:85:Control.fir@5.4]
  output        io_ctrl_Branch_Src, // @[control.py:85:Control.fir@5.4]
  output        io_ctrl_Mem_Read, // @[control.py:85:Control.fir@5.4]
  output        io_ctrl_Mem_Write, // @[control.py:85:Control.fir@5.4]
  output [1:0]  io_ctrl_Data_Size, // @[control.py:85:Control.fir@5.4]
  output        io_ctrl_Load_Type, // @[control.py:85:Control.fir@5.4]
  output [2:0]  io_ctrl_Mem_to_Reg, // @[control.py:85:Control.fir@5.4]
  output        io_ctrl_Jump_Type // @[control.py:85:Control.fir@5.4]
);
  wire [31:0] _T_19; // @[listlookup.py:52:Control.fir@7.4]
  wire  _T_20; // @[listlookup.py:52:Control.fir@8.4]
  wire  _T_22; // @[listlookup.py:52:Control.fir@10.4]
  wire  _T_24; // @[listlookup.py:52:Control.fir@12.4]
  wire  _T_26; // @[listlookup.py:52:Control.fir@14.4]
  wire  _T_28; // @[listlookup.py:52:Control.fir@16.4]
  wire [31:0] _T_29; // @[listlookup.py:52:Control.fir@17.4]
  wire  _T_30; // @[listlookup.py:52:Control.fir@18.4]
  wire  _T_32; // @[listlookup.py:52:Control.fir@20.4]
  wire  _T_34; // @[listlookup.py:52:Control.fir@22.4]
  wire  _T_36; // @[listlookup.py:52:Control.fir@24.4]
  wire  _T_38; // @[listlookup.py:52:Control.fir@26.4]
  wire  _T_40; // @[listlookup.py:52:Control.fir@28.4]
  wire  _T_42; // @[listlookup.py:52:Control.fir@30.4]
  wire  _T_44; // @[listlookup.py:52:Control.fir@32.4]
  wire  _T_46; // @[listlookup.py:52:Control.fir@34.4]
  wire  _T_48; // @[listlookup.py:52:Control.fir@36.4]
  wire  _T_50; // @[listlookup.py:52:Control.fir@38.4]
  wire  _T_52; // @[listlookup.py:52:Control.fir@40.4]
  wire  _T_54; // @[listlookup.py:52:Control.fir@42.4]
  wire  _T_56; // @[listlookup.py:52:Control.fir@44.4]
  wire  _T_58; // @[listlookup.py:52:Control.fir@46.4]
  wire  _T_60; // @[listlookup.py:52:Control.fir@48.4]
  wire  _T_62; // @[listlookup.py:52:Control.fir@50.4]
  wire  _T_64; // @[listlookup.py:52:Control.fir@52.4]
  wire  _T_66; // @[listlookup.py:52:Control.fir@54.4]
  wire  _T_68; // @[listlookup.py:52:Control.fir@56.4]
  wire  _T_70; // @[listlookup.py:52:Control.fir@58.4]
  wire  _T_72; // @[listlookup.py:52:Control.fir@60.4]
  wire  _T_74; // @[listlookup.py:52:Control.fir@62.4]
  wire  _T_76; // @[listlookup.py:52:Control.fir@64.4]
  wire  _T_78; // @[listlookup.py:52:Control.fir@66.4]
  wire  _T_80; // @[listlookup.py:52:Control.fir@68.4]
  wire  _T_82; // @[listlookup.py:52:Control.fir@70.4]
  wire  _T_84; // @[listlookup.py:52:Control.fir@72.4]
  wire [31:0] _T_85; // @[listlookup.py:52:Control.fir@73.4]
  wire  _T_86; // @[listlookup.py:52:Control.fir@74.4]
  wire  _T_88; // @[listlookup.py:52:Control.fir@76.4]
  wire  _T_90; // @[listlookup.py:52:Control.fir@78.4]
  wire  _T_92; // @[listlookup.py:52:Control.fir@80.4]
  wire  _T_97; // @[control.py:95:Control.fir@85.4]
  wire  _T_98; // @[control.py:95:Control.fir@86.4]
  wire  _T_99; // @[control.py:95:Control.fir@87.4]
  wire  _T_100; // @[control.py:95:Control.fir@88.4]
  wire  _T_101; // @[control.py:95:Control.fir@89.4]
  wire  _T_102; // @[control.py:95:Control.fir@90.4]
  wire  _T_103; // @[control.py:95:Control.fir@91.4]
  wire  _T_104; // @[control.py:95:Control.fir@92.4]
  wire  _T_105; // @[control.py:95:Control.fir@93.4]
  wire  _T_106; // @[control.py:95:Control.fir@94.4]
  wire  _T_107; // @[control.py:95:Control.fir@95.4]
  wire  _T_108; // @[control.py:95:Control.fir@96.4]
  wire  _T_109; // @[control.py:95:Control.fir@97.4]
  wire  _T_110; // @[control.py:95:Control.fir@98.4]
  wire  _T_111; // @[control.py:95:Control.fir@99.4]
  wire  _T_112; // @[control.py:95:Control.fir@100.4]
  wire  _T_113; // @[control.py:95:Control.fir@101.4]
  wire  _T_114; // @[control.py:95:Control.fir@102.4]
  wire  _T_115; // @[control.py:95:Control.fir@103.4]
  wire  _T_116; // @[control.py:95:Control.fir@104.4]
  wire  _T_117; // @[control.py:95:Control.fir@105.4]
  wire  _T_118; // @[control.py:95:Control.fir@106.4]
  wire  _T_119; // @[control.py:95:Control.fir@107.4]
  wire  _T_120; // @[control.py:95:Control.fir@108.4]
  wire  _T_121; // @[control.py:95:Control.fir@109.4]
  wire  _T_122; // @[control.py:95:Control.fir@110.4]
  wire  _T_123; // @[control.py:95:Control.fir@111.4]
  wire  _T_124; // @[control.py:95:Control.fir@112.4]
  wire  _T_125; // @[control.py:95:Control.fir@113.4]
  wire  _T_126; // @[control.py:95:Control.fir@114.4]
  wire  _T_127; // @[control.py:95:Control.fir@115.4]
  wire  _T_128; // @[control.py:95:Control.fir@116.4]
  wire  _T_129; // @[control.py:95:Control.fir@117.4]
  wire  _T_130; // @[control.py:95:Control.fir@118.4]
  wire  _T_131; // @[control.py:95:Control.fir@119.4]
  wire [2:0] _T_134; // @[control.py:95:Control.fir@122.4]
  wire [2:0] _T_135; // @[control.py:95:Control.fir@123.4]
  wire [2:0] _T_136; // @[control.py:95:Control.fir@124.4]
  wire [2:0] _T_137; // @[control.py:95:Control.fir@125.4]
  wire [2:0] _T_138; // @[control.py:95:Control.fir@126.4]
  wire [2:0] _T_139; // @[control.py:95:Control.fir@127.4]
  wire [2:0] _T_140; // @[control.py:95:Control.fir@128.4]
  wire [2:0] _T_141; // @[control.py:95:Control.fir@129.4]
  wire [2:0] _T_142; // @[control.py:95:Control.fir@130.4]
  wire [2:0] _T_143; // @[control.py:95:Control.fir@131.4]
  wire [2:0] _T_144; // @[control.py:95:Control.fir@132.4]
  wire [2:0] _T_145; // @[control.py:95:Control.fir@133.4]
  wire [2:0] _T_146; // @[control.py:95:Control.fir@134.4]
  wire [2:0] _T_147; // @[control.py:95:Control.fir@135.4]
  wire [2:0] _T_148; // @[control.py:95:Control.fir@136.4]
  wire [2:0] _T_149; // @[control.py:95:Control.fir@137.4]
  wire [2:0] _T_150; // @[control.py:95:Control.fir@138.4]
  wire [2:0] _T_151; // @[control.py:95:Control.fir@139.4]
  wire [2:0] _T_152; // @[control.py:95:Control.fir@140.4]
  wire [2:0] _T_153; // @[control.py:95:Control.fir@141.4]
  wire [2:0] _T_154; // @[control.py:95:Control.fir@142.4]
  wire [2:0] _T_155; // @[control.py:95:Control.fir@143.4]
  wire [2:0] _T_156; // @[control.py:95:Control.fir@144.4]
  wire [2:0] _T_157; // @[control.py:95:Control.fir@145.4]
  wire [2:0] _T_158; // @[control.py:95:Control.fir@146.4]
  wire [2:0] _T_159; // @[control.py:95:Control.fir@147.4]
  wire [2:0] _T_160; // @[control.py:95:Control.fir@148.4]
  wire [2:0] _T_161; // @[control.py:95:Control.fir@149.4]
  wire [2:0] _T_162; // @[control.py:95:Control.fir@150.4]
  wire [2:0] _T_163; // @[control.py:95:Control.fir@151.4]
  wire [2:0] _T_164; // @[control.py:95:Control.fir@152.4]
  wire [2:0] _T_165; // @[control.py:95:Control.fir@153.4]
  wire [2:0] _T_166; // @[control.py:95:Control.fir@154.4]
  wire [2:0] _T_167; // @[control.py:95:Control.fir@155.4]
  wire [2:0] _T_168; // @[control.py:95:Control.fir@156.4]
  wire [2:0] _T_169; // @[control.py:95:Control.fir@157.4]
  wire  _T_183; // @[control.py:95:Control.fir@171.4]
  wire  _T_184; // @[control.py:95:Control.fir@172.4]
  wire  _T_185; // @[control.py:95:Control.fir@173.4]
  wire  _T_186; // @[control.py:95:Control.fir@174.4]
  wire  _T_187; // @[control.py:95:Control.fir@175.4]
  wire  _T_188; // @[control.py:95:Control.fir@176.4]
  wire  _T_189; // @[control.py:95:Control.fir@177.4]
  wire  _T_190; // @[control.py:95:Control.fir@178.4]
  wire  _T_191; // @[control.py:95:Control.fir@179.4]
  wire  _T_192; // @[control.py:95:Control.fir@180.4]
  wire  _T_193; // @[control.py:95:Control.fir@181.4]
  wire  _T_194; // @[control.py:95:Control.fir@182.4]
  wire  _T_195; // @[control.py:95:Control.fir@183.4]
  wire  _T_196; // @[control.py:95:Control.fir@184.4]
  wire  _T_197; // @[control.py:95:Control.fir@185.4]
  wire  _T_198; // @[control.py:95:Control.fir@186.4]
  wire  _T_199; // @[control.py:95:Control.fir@187.4]
  wire  _T_200; // @[control.py:95:Control.fir@188.4]
  wire  _T_201; // @[control.py:95:Control.fir@189.4]
  wire  _T_202; // @[control.py:95:Control.fir@190.4]
  wire  _T_203; // @[control.py:95:Control.fir@191.4]
  wire  _T_204; // @[control.py:95:Control.fir@192.4]
  wire  _T_205; // @[control.py:95:Control.fir@193.4]
  wire  _T_206; // @[control.py:95:Control.fir@194.4]
  wire  _T_207; // @[control.py:95:Control.fir@195.4]
  wire [4:0] _T_210; // @[control.py:95:Control.fir@198.4]
  wire [4:0] _T_211; // @[control.py:95:Control.fir@199.4]
  wire [4:0] _T_212; // @[control.py:95:Control.fir@200.4]
  wire [4:0] _T_213; // @[control.py:95:Control.fir@201.4]
  wire [4:0] _T_214; // @[control.py:95:Control.fir@202.4]
  wire [4:0] _T_215; // @[control.py:95:Control.fir@203.4]
  wire [4:0] _T_216; // @[control.py:95:Control.fir@204.4]
  wire [4:0] _T_217; // @[control.py:95:Control.fir@205.4]
  wire [4:0] _T_218; // @[control.py:95:Control.fir@206.4]
  wire [4:0] _T_219; // @[control.py:95:Control.fir@207.4]
  wire [4:0] _T_220; // @[control.py:95:Control.fir@208.4]
  wire [4:0] _T_221; // @[control.py:95:Control.fir@209.4]
  wire [4:0] _T_222; // @[control.py:95:Control.fir@210.4]
  wire [4:0] _T_223; // @[control.py:95:Control.fir@211.4]
  wire [4:0] _T_224; // @[control.py:95:Control.fir@212.4]
  wire [4:0] _T_225; // @[control.py:95:Control.fir@213.4]
  wire [4:0] _T_226; // @[control.py:95:Control.fir@214.4]
  wire [4:0] _T_227; // @[control.py:95:Control.fir@215.4]
  wire [4:0] _T_228; // @[control.py:95:Control.fir@216.4]
  wire [4:0] _T_229; // @[control.py:95:Control.fir@217.4]
  wire [4:0] _T_230; // @[control.py:95:Control.fir@218.4]
  wire [4:0] _T_231; // @[control.py:95:Control.fir@219.4]
  wire [4:0] _T_232; // @[control.py:95:Control.fir@220.4]
  wire [4:0] _T_233; // @[control.py:95:Control.fir@221.4]
  wire [4:0] _T_234; // @[control.py:95:Control.fir@222.4]
  wire [4:0] _T_235; // @[control.py:95:Control.fir@223.4]
  wire [4:0] _T_236; // @[control.py:95:Control.fir@224.4]
  wire [4:0] _T_237; // @[control.py:95:Control.fir@225.4]
  wire [4:0] _T_238; // @[control.py:95:Control.fir@226.4]
  wire [4:0] _T_239; // @[control.py:95:Control.fir@227.4]
  wire [4:0] _T_240; // @[control.py:95:Control.fir@228.4]
  wire [4:0] _T_241; // @[control.py:95:Control.fir@229.4]
  wire [4:0] _T_242; // @[control.py:95:Control.fir@230.4]
  wire [4:0] _T_243; // @[control.py:95:Control.fir@231.4]
  wire [4:0] _T_244; // @[control.py:95:Control.fir@232.4]
  wire [4:0] _T_245; // @[control.py:95:Control.fir@233.4]
  wire  _T_251; // @[control.py:95:Control.fir@239.4]
  wire  _T_252; // @[control.py:95:Control.fir@240.4]
  wire  _T_253; // @[control.py:95:Control.fir@241.4]
  wire  _T_254; // @[control.py:95:Control.fir@242.4]
  wire  _T_255; // @[control.py:95:Control.fir@243.4]
  wire  _T_256; // @[control.py:95:Control.fir@244.4]
  wire  _T_257; // @[control.py:95:Control.fir@245.4]
  wire  _T_258; // @[control.py:95:Control.fir@246.4]
  wire  _T_259; // @[control.py:95:Control.fir@247.4]
  wire  _T_260; // @[control.py:95:Control.fir@248.4]
  wire  _T_261; // @[control.py:95:Control.fir@249.4]
  wire  _T_262; // @[control.py:95:Control.fir@250.4]
  wire  _T_263; // @[control.py:95:Control.fir@251.4]
  wire  _T_264; // @[control.py:95:Control.fir@252.4]
  wire  _T_265; // @[control.py:95:Control.fir@253.4]
  wire  _T_266; // @[control.py:95:Control.fir@254.4]
  wire  _T_267; // @[control.py:95:Control.fir@255.4]
  wire  _T_268; // @[control.py:95:Control.fir@256.4]
  wire  _T_269; // @[control.py:95:Control.fir@257.4]
  wire  _T_270; // @[control.py:95:Control.fir@258.4]
  wire  _T_271; // @[control.py:95:Control.fir@259.4]
  wire  _T_272; // @[control.py:95:Control.fir@260.4]
  wire  _T_273; // @[control.py:95:Control.fir@261.4]
  wire  _T_274; // @[control.py:95:Control.fir@262.4]
  wire  _T_275; // @[control.py:95:Control.fir@263.4]
  wire  _T_276; // @[control.py:95:Control.fir@264.4]
  wire  _T_277; // @[control.py:95:Control.fir@265.4]
  wire  _T_278; // @[control.py:95:Control.fir@266.4]
  wire  _T_279; // @[control.py:95:Control.fir@267.4]
  wire  _T_280; // @[control.py:95:Control.fir@268.4]
  wire  _T_281; // @[control.py:95:Control.fir@269.4]
  wire  _T_282; // @[control.py:95:Control.fir@270.4]
  wire  _T_283; // @[control.py:95:Control.fir@271.4]
  wire  _T_289; // @[control.py:95:Control.fir@277.4]
  wire  _T_290; // @[control.py:95:Control.fir@278.4]
  wire  _T_291; // @[control.py:95:Control.fir@279.4]
  wire  _T_292; // @[control.py:95:Control.fir@280.4]
  wire  _T_293; // @[control.py:95:Control.fir@281.4]
  wire  _T_294; // @[control.py:95:Control.fir@282.4]
  wire  _T_295; // @[control.py:95:Control.fir@283.4]
  wire  _T_296; // @[control.py:95:Control.fir@284.4]
  wire  _T_297; // @[control.py:95:Control.fir@285.4]
  wire  _T_298; // @[control.py:95:Control.fir@286.4]
  wire  _T_299; // @[control.py:95:Control.fir@287.4]
  wire  _T_300; // @[control.py:95:Control.fir@288.4]
  wire  _T_301; // @[control.py:95:Control.fir@289.4]
  wire  _T_302; // @[control.py:95:Control.fir@290.4]
  wire  _T_303; // @[control.py:95:Control.fir@291.4]
  wire  _T_304; // @[control.py:95:Control.fir@292.4]
  wire  _T_305; // @[control.py:95:Control.fir@293.4]
  wire  _T_306; // @[control.py:95:Control.fir@294.4]
  wire  _T_307; // @[control.py:95:Control.fir@295.4]
  wire  _T_308; // @[control.py:95:Control.fir@296.4]
  wire  _T_309; // @[control.py:95:Control.fir@297.4]
  wire  _T_310; // @[control.py:95:Control.fir@298.4]
  wire  _T_311; // @[control.py:95:Control.fir@299.4]
  wire  _T_312; // @[control.py:95:Control.fir@300.4]
  wire  _T_313; // @[control.py:95:Control.fir@301.4]
  wire  _T_314; // @[control.py:95:Control.fir@302.4]
  wire  _T_315; // @[control.py:95:Control.fir@303.4]
  wire  _T_316; // @[control.py:95:Control.fir@304.4]
  wire  _T_317; // @[control.py:95:Control.fir@305.4]
  wire  _T_318; // @[control.py:95:Control.fir@306.4]
  wire  _T_319; // @[control.py:95:Control.fir@307.4]
  wire  _T_320; // @[control.py:95:Control.fir@308.4]
  wire  _T_321; // @[control.py:95:Control.fir@309.4]
  wire  _T_338; // @[control.py:95:Control.fir@326.4]
  wire  _T_339; // @[control.py:95:Control.fir@327.4]
  wire  _T_340; // @[control.py:95:Control.fir@328.4]
  wire  _T_341; // @[control.py:95:Control.fir@329.4]
  wire  _T_342; // @[control.py:95:Control.fir@330.4]
  wire  _T_343; // @[control.py:95:Control.fir@331.4]
  wire  _T_344; // @[control.py:95:Control.fir@332.4]
  wire  _T_345; // @[control.py:95:Control.fir@333.4]
  wire  _T_346; // @[control.py:95:Control.fir@334.4]
  wire  _T_347; // @[control.py:95:Control.fir@335.4]
  wire  _T_348; // @[control.py:95:Control.fir@336.4]
  wire  _T_349; // @[control.py:95:Control.fir@337.4]
  wire  _T_350; // @[control.py:95:Control.fir@338.4]
  wire  _T_351; // @[control.py:95:Control.fir@339.4]
  wire  _T_352; // @[control.py:95:Control.fir@340.4]
  wire  _T_353; // @[control.py:95:Control.fir@341.4]
  wire  _T_354; // @[control.py:95:Control.fir@342.4]
  wire  _T_355; // @[control.py:95:Control.fir@343.4]
  wire  _T_356; // @[control.py:95:Control.fir@344.4]
  wire  _T_357; // @[control.py:95:Control.fir@345.4]
  wire  _T_358; // @[control.py:95:Control.fir@346.4]
  wire  _T_359; // @[control.py:95:Control.fir@347.4]
  wire  _T_375; // @[control.py:95:Control.fir@363.4]
  wire  _T_376; // @[control.py:95:Control.fir@364.4]
  wire  _T_377; // @[control.py:95:Control.fir@365.4]
  wire  _T_378; // @[control.py:95:Control.fir@366.4]
  wire  _T_379; // @[control.py:95:Control.fir@367.4]
  wire  _T_380; // @[control.py:95:Control.fir@368.4]
  wire  _T_381; // @[control.py:95:Control.fir@369.4]
  wire  _T_382; // @[control.py:95:Control.fir@370.4]
  wire  _T_383; // @[control.py:95:Control.fir@371.4]
  wire  _T_384; // @[control.py:95:Control.fir@372.4]
  wire  _T_385; // @[control.py:95:Control.fir@373.4]
  wire  _T_386; // @[control.py:95:Control.fir@374.4]
  wire  _T_387; // @[control.py:95:Control.fir@375.4]
  wire  _T_388; // @[control.py:95:Control.fir@376.4]
  wire  _T_389; // @[control.py:95:Control.fir@377.4]
  wire  _T_390; // @[control.py:95:Control.fir@378.4]
  wire  _T_391; // @[control.py:95:Control.fir@379.4]
  wire  _T_392; // @[control.py:95:Control.fir@380.4]
  wire  _T_393; // @[control.py:95:Control.fir@381.4]
  wire  _T_394; // @[control.py:95:Control.fir@382.4]
  wire  _T_395; // @[control.py:95:Control.fir@383.4]
  wire  _T_396; // @[control.py:95:Control.fir@384.4]
  wire  _T_397; // @[control.py:95:Control.fir@385.4]
  wire [1:0] _T_410; // @[control.py:95:Control.fir@398.4]
  wire [1:0] _T_411; // @[control.py:95:Control.fir@399.4]
  wire [1:0] _T_412; // @[control.py:95:Control.fir@400.4]
  wire [1:0] _T_413; // @[control.py:95:Control.fir@401.4]
  wire [1:0] _T_414; // @[control.py:95:Control.fir@402.4]
  wire [1:0] _T_415; // @[control.py:95:Control.fir@403.4]
  wire [1:0] _T_416; // @[control.py:95:Control.fir@404.4]
  wire [1:0] _T_417; // @[control.py:95:Control.fir@405.4]
  wire [1:0] _T_418; // @[control.py:95:Control.fir@406.4]
  wire [1:0] _T_419; // @[control.py:95:Control.fir@407.4]
  wire [1:0] _T_420; // @[control.py:95:Control.fir@408.4]
  wire [1:0] _T_421; // @[control.py:95:Control.fir@409.4]
  wire [1:0] _T_422; // @[control.py:95:Control.fir@410.4]
  wire [1:0] _T_423; // @[control.py:95:Control.fir@411.4]
  wire [1:0] _T_424; // @[control.py:95:Control.fir@412.4]
  wire [1:0] _T_425; // @[control.py:95:Control.fir@413.4]
  wire [1:0] _T_426; // @[control.py:95:Control.fir@414.4]
  wire [1:0] _T_427; // @[control.py:95:Control.fir@415.4]
  wire [1:0] _T_428; // @[control.py:95:Control.fir@416.4]
  wire [1:0] _T_429; // @[control.py:95:Control.fir@417.4]
  wire [1:0] _T_430; // @[control.py:95:Control.fir@418.4]
  wire [1:0] _T_431; // @[control.py:95:Control.fir@419.4]
  wire [1:0] _T_432; // @[control.py:95:Control.fir@420.4]
  wire [1:0] _T_433; // @[control.py:95:Control.fir@421.4]
  wire [1:0] _T_434; // @[control.py:95:Control.fir@422.4]
  wire [1:0] _T_435; // @[control.py:95:Control.fir@423.4]
  wire  _T_453; // @[control.py:95:Control.fir@441.4]
  wire  _T_454; // @[control.py:95:Control.fir@442.4]
  wire  _T_455; // @[control.py:95:Control.fir@443.4]
  wire  _T_456; // @[control.py:95:Control.fir@444.4]
  wire  _T_457; // @[control.py:95:Control.fir@445.4]
  wire  _T_458; // @[control.py:95:Control.fir@446.4]
  wire  _T_459; // @[control.py:95:Control.fir@447.4]
  wire  _T_460; // @[control.py:95:Control.fir@448.4]
  wire  _T_461; // @[control.py:95:Control.fir@449.4]
  wire  _T_462; // @[control.py:95:Control.fir@450.4]
  wire  _T_463; // @[control.py:95:Control.fir@451.4]
  wire  _T_464; // @[control.py:95:Control.fir@452.4]
  wire  _T_465; // @[control.py:95:Control.fir@453.4]
  wire  _T_466; // @[control.py:95:Control.fir@454.4]
  wire  _T_467; // @[control.py:95:Control.fir@455.4]
  wire  _T_468; // @[control.py:95:Control.fir@456.4]
  wire  _T_469; // @[control.py:95:Control.fir@457.4]
  wire  _T_470; // @[control.py:95:Control.fir@458.4]
  wire  _T_471; // @[control.py:95:Control.fir@459.4]
  wire  _T_472; // @[control.py:95:Control.fir@460.4]
  wire  _T_473; // @[control.py:95:Control.fir@461.4]
  wire [2:0] _T_476; // @[control.py:95:Control.fir@464.4]
  wire [2:0] _T_477; // @[control.py:95:Control.fir@465.4]
  wire [2:0] _T_478; // @[control.py:95:Control.fir@466.4]
  wire [2:0] _T_479; // @[control.py:95:Control.fir@467.4]
  wire [2:0] _T_480; // @[control.py:95:Control.fir@468.4]
  wire [2:0] _T_481; // @[control.py:95:Control.fir@469.4]
  wire [2:0] _T_482; // @[control.py:95:Control.fir@470.4]
  wire [2:0] _T_483; // @[control.py:95:Control.fir@471.4]
  wire [2:0] _T_484; // @[control.py:95:Control.fir@472.4]
  wire [2:0] _T_485; // @[control.py:95:Control.fir@473.4]
  wire [2:0] _T_486; // @[control.py:95:Control.fir@474.4]
  wire [2:0] _T_487; // @[control.py:95:Control.fir@475.4]
  wire [2:0] _T_488; // @[control.py:95:Control.fir@476.4]
  wire [2:0] _T_489; // @[control.py:95:Control.fir@477.4]
  wire [2:0] _T_490; // @[control.py:95:Control.fir@478.4]
  wire [2:0] _T_491; // @[control.py:95:Control.fir@479.4]
  wire [2:0] _T_492; // @[control.py:95:Control.fir@480.4]
  wire [2:0] _T_493; // @[control.py:95:Control.fir@481.4]
  wire [2:0] _T_494; // @[control.py:95:Control.fir@482.4]
  wire [2:0] _T_495; // @[control.py:95:Control.fir@483.4]
  wire [2:0] _T_496; // @[control.py:95:Control.fir@484.4]
  wire [2:0] _T_497; // @[control.py:95:Control.fir@485.4]
  wire [2:0] _T_498; // @[control.py:95:Control.fir@486.4]
  wire [2:0] _T_499; // @[control.py:95:Control.fir@487.4]
  wire [2:0] _T_500; // @[control.py:95:Control.fir@488.4]
  wire [2:0] _T_501; // @[control.py:95:Control.fir@489.4]
  wire [2:0] _T_502; // @[control.py:95:Control.fir@490.4]
  wire [2:0] _T_503; // @[control.py:95:Control.fir@491.4]
  wire [2:0] _T_504; // @[control.py:95:Control.fir@492.4]
  wire [2:0] _T_505; // @[control.py:95:Control.fir@493.4]
  wire [2:0] _T_506; // @[control.py:95:Control.fir@494.4]
  wire [2:0] _T_507; // @[control.py:95:Control.fir@495.4]
  wire [2:0] _T_508; // @[control.py:95:Control.fir@496.4]
  wire [2:0] _T_509; // @[control.py:95:Control.fir@497.4]
  wire [2:0] _T_510; // @[control.py:95:Control.fir@498.4]
  wire [2:0] _T_511; // @[control.py:95:Control.fir@499.4]
  wire  _T_518; // @[control.py:95:Control.fir@506.4]
  wire  _T_519; // @[control.py:95:Control.fir@507.4]
  wire  _T_520; // @[control.py:95:Control.fir@508.4]
  wire  _T_521; // @[control.py:95:Control.fir@509.4]
  wire  _T_522; // @[control.py:95:Control.fir@510.4]
  wire  _T_523; // @[control.py:95:Control.fir@511.4]
  wire  _T_524; // @[control.py:95:Control.fir@512.4]
  wire  _T_525; // @[control.py:95:Control.fir@513.4]
  wire  _T_526; // @[control.py:95:Control.fir@514.4]
  wire  _T_527; // @[control.py:95:Control.fir@515.4]
  wire  _T_528; // @[control.py:95:Control.fir@516.4]
  wire  _T_529; // @[control.py:95:Control.fir@517.4]
  wire  _T_530; // @[control.py:95:Control.fir@518.4]
  wire  _T_531; // @[control.py:95:Control.fir@519.4]
  wire  _T_532; // @[control.py:95:Control.fir@520.4]
  wire  _T_533; // @[control.py:95:Control.fir@521.4]
  wire  _T_534; // @[control.py:95:Control.fir@522.4]
  wire  _T_535; // @[control.py:95:Control.fir@523.4]
  wire  _T_536; // @[control.py:95:Control.fir@524.4]
  wire  _T_537; // @[control.py:95:Control.fir@525.4]
  wire  _T_538; // @[control.py:95:Control.fir@526.4]
  wire  _T_539; // @[control.py:95:Control.fir@527.4]
  wire  _T_540; // @[control.py:95:Control.fir@528.4]
  wire  _T_541; // @[control.py:95:Control.fir@529.4]
  wire  _T_542; // @[control.py:95:Control.fir@530.4]
  wire  _T_543; // @[control.py:95:Control.fir@531.4]
  wire  _T_544; // @[control.py:95:Control.fir@532.4]
  wire  _T_545; // @[control.py:95:Control.fir@533.4]
  wire  _T_546; // @[control.py:95:Control.fir@534.4]
  wire  _T_547; // @[control.py:95:Control.fir@535.4]
  wire  _T_548; // @[control.py:95:Control.fir@536.4]
  wire  _T_549; // @[control.py:95:Control.fir@537.4]
  assign _T_19 = io_inst & 32'hfe00707f; // @[listlookup.py:52:Control.fir@7.4]
  assign _T_20 = _T_19 == 32'h33; // @[listlookup.py:52:Control.fir@8.4]
  assign _T_22 = _T_19 == 32'h40000033; // @[listlookup.py:52:Control.fir@10.4]
  assign _T_24 = _T_19 == 32'h7033; // @[listlookup.py:52:Control.fir@12.4]
  assign _T_26 = _T_19 == 32'h6033; // @[listlookup.py:52:Control.fir@14.4]
  assign _T_28 = _T_19 == 32'h4033; // @[listlookup.py:52:Control.fir@16.4]
  assign _T_29 = io_inst & 32'h707f; // @[listlookup.py:52:Control.fir@17.4]
  assign _T_30 = _T_29 == 32'h13; // @[listlookup.py:52:Control.fir@18.4]
  assign _T_32 = _T_29 == 32'h7013; // @[listlookup.py:52:Control.fir@20.4]
  assign _T_34 = _T_29 == 32'h6013; // @[listlookup.py:52:Control.fir@22.4]
  assign _T_36 = _T_29 == 32'h4013; // @[listlookup.py:52:Control.fir@24.4]
  assign _T_38 = _T_19 == 32'h1033; // @[listlookup.py:52:Control.fir@26.4]
  assign _T_40 = _T_19 == 32'h5033; // @[listlookup.py:52:Control.fir@28.4]
  assign _T_42 = _T_19 == 32'h40005033; // @[listlookup.py:52:Control.fir@30.4]
  assign _T_44 = _T_19 == 32'h1013; // @[listlookup.py:52:Control.fir@32.4]
  assign _T_46 = _T_19 == 32'h5013; // @[listlookup.py:52:Control.fir@34.4]
  assign _T_48 = _T_19 == 32'h40005013; // @[listlookup.py:52:Control.fir@36.4]
  assign _T_50 = _T_19 == 32'h2033; // @[listlookup.py:52:Control.fir@38.4]
  assign _T_52 = _T_19 == 32'h3033; // @[listlookup.py:52:Control.fir@40.4]
  assign _T_54 = _T_29 == 32'h2013; // @[listlookup.py:52:Control.fir@42.4]
  assign _T_56 = _T_29 == 32'h3013; // @[listlookup.py:52:Control.fir@44.4]
  assign _T_58 = _T_29 == 32'h2003; // @[listlookup.py:52:Control.fir@46.4]
  assign _T_60 = _T_29 == 32'h1003; // @[listlookup.py:52:Control.fir@48.4]
  assign _T_62 = _T_29 == 32'h3; // @[listlookup.py:52:Control.fir@50.4]
  assign _T_64 = _T_29 == 32'h5003; // @[listlookup.py:52:Control.fir@52.4]
  assign _T_66 = _T_29 == 32'h4003; // @[listlookup.py:52:Control.fir@54.4]
  assign _T_68 = _T_29 == 32'h2023; // @[listlookup.py:52:Control.fir@56.4]
  assign _T_70 = _T_29 == 32'h1023; // @[listlookup.py:52:Control.fir@58.4]
  assign _T_72 = _T_29 == 32'h23; // @[listlookup.py:52:Control.fir@60.4]
  assign _T_74 = _T_29 == 32'h63; // @[listlookup.py:52:Control.fir@62.4]
  assign _T_76 = _T_29 == 32'h1063; // @[listlookup.py:52:Control.fir@64.4]
  assign _T_78 = _T_29 == 32'h4063; // @[listlookup.py:52:Control.fir@66.4]
  assign _T_80 = _T_29 == 32'h5063; // @[listlookup.py:52:Control.fir@68.4]
  assign _T_82 = _T_29 == 32'h6063; // @[listlookup.py:52:Control.fir@70.4]
  assign _T_84 = _T_29 == 32'h7063; // @[listlookup.py:52:Control.fir@72.4]
  assign _T_85 = io_inst & 32'h7f; // @[listlookup.py:52:Control.fir@73.4]
  assign _T_86 = _T_85 == 32'h6f; // @[listlookup.py:52:Control.fir@74.4]
  assign _T_88 = _T_29 == 32'h67; // @[listlookup.py:52:Control.fir@76.4]
  assign _T_90 = _T_85 == 32'h37; // @[listlookup.py:52:Control.fir@78.4]
  assign _T_92 = _T_85 == 32'h17; // @[listlookup.py:52:Control.fir@80.4]
  assign _T_97 = _T_90 ? 1'h1 : _T_92; // @[control.py:95:Control.fir@85.4]
  assign _T_98 = _T_88 ? 1'h1 : _T_97; // @[control.py:95:Control.fir@86.4]
  assign _T_99 = _T_86 ? 1'h1 : _T_98; // @[control.py:95:Control.fir@87.4]
  assign _T_100 = _T_84 ? 1'h0 : _T_99; // @[control.py:95:Control.fir@88.4]
  assign _T_101 = _T_82 ? 1'h0 : _T_100; // @[control.py:95:Control.fir@89.4]
  assign _T_102 = _T_80 ? 1'h0 : _T_101; // @[control.py:95:Control.fir@90.4]
  assign _T_103 = _T_78 ? 1'h0 : _T_102; // @[control.py:95:Control.fir@91.4]
  assign _T_104 = _T_76 ? 1'h0 : _T_103; // @[control.py:95:Control.fir@92.4]
  assign _T_105 = _T_74 ? 1'h0 : _T_104; // @[control.py:95:Control.fir@93.4]
  assign _T_106 = _T_72 ? 1'h0 : _T_105; // @[control.py:95:Control.fir@94.4]
  assign _T_107 = _T_70 ? 1'h0 : _T_106; // @[control.py:95:Control.fir@95.4]
  assign _T_108 = _T_68 ? 1'h0 : _T_107; // @[control.py:95:Control.fir@96.4]
  assign _T_109 = _T_66 ? 1'h1 : _T_108; // @[control.py:95:Control.fir@97.4]
  assign _T_110 = _T_64 ? 1'h1 : _T_109; // @[control.py:95:Control.fir@98.4]
  assign _T_111 = _T_62 ? 1'h1 : _T_110; // @[control.py:95:Control.fir@99.4]
  assign _T_112 = _T_60 ? 1'h1 : _T_111; // @[control.py:95:Control.fir@100.4]
  assign _T_113 = _T_58 ? 1'h1 : _T_112; // @[control.py:95:Control.fir@101.4]
  assign _T_114 = _T_56 ? 1'h1 : _T_113; // @[control.py:95:Control.fir@102.4]
  assign _T_115 = _T_54 ? 1'h1 : _T_114; // @[control.py:95:Control.fir@103.4]
  assign _T_116 = _T_52 ? 1'h1 : _T_115; // @[control.py:95:Control.fir@104.4]
  assign _T_117 = _T_50 ? 1'h1 : _T_116; // @[control.py:95:Control.fir@105.4]
  assign _T_118 = _T_48 ? 1'h1 : _T_117; // @[control.py:95:Control.fir@106.4]
  assign _T_119 = _T_46 ? 1'h1 : _T_118; // @[control.py:95:Control.fir@107.4]
  assign _T_120 = _T_44 ? 1'h1 : _T_119; // @[control.py:95:Control.fir@108.4]
  assign _T_121 = _T_42 ? 1'h1 : _T_120; // @[control.py:95:Control.fir@109.4]
  assign _T_122 = _T_40 ? 1'h1 : _T_121; // @[control.py:95:Control.fir@110.4]
  assign _T_123 = _T_38 ? 1'h1 : _T_122; // @[control.py:95:Control.fir@111.4]
  assign _T_124 = _T_36 ? 1'h1 : _T_123; // @[control.py:95:Control.fir@112.4]
  assign _T_125 = _T_34 ? 1'h1 : _T_124; // @[control.py:95:Control.fir@113.4]
  assign _T_126 = _T_32 ? 1'h1 : _T_125; // @[control.py:95:Control.fir@114.4]
  assign _T_127 = _T_30 ? 1'h1 : _T_126; // @[control.py:95:Control.fir@115.4]
  assign _T_128 = _T_28 ? 1'h1 : _T_127; // @[control.py:95:Control.fir@116.4]
  assign _T_129 = _T_26 ? 1'h1 : _T_128; // @[control.py:95:Control.fir@117.4]
  assign _T_130 = _T_24 ? 1'h1 : _T_129; // @[control.py:95:Control.fir@118.4]
  assign _T_131 = _T_22 ? 1'h1 : _T_130; // @[control.py:95:Control.fir@119.4]
  assign _T_134 = _T_92 ? 3'h5 : 3'h0; // @[control.py:95:Control.fir@122.4]
  assign _T_135 = _T_90 ? 3'h5 : _T_134; // @[control.py:95:Control.fir@123.4]
  assign _T_136 = _T_88 ? 3'h2 : _T_135; // @[control.py:95:Control.fir@124.4]
  assign _T_137 = _T_86 ? 3'h6 : _T_136; // @[control.py:95:Control.fir@125.4]
  assign _T_138 = _T_84 ? 3'h4 : _T_137; // @[control.py:95:Control.fir@126.4]
  assign _T_139 = _T_82 ? 3'h4 : _T_138; // @[control.py:95:Control.fir@127.4]
  assign _T_140 = _T_80 ? 3'h4 : _T_139; // @[control.py:95:Control.fir@128.4]
  assign _T_141 = _T_78 ? 3'h4 : _T_140; // @[control.py:95:Control.fir@129.4]
  assign _T_142 = _T_76 ? 3'h4 : _T_141; // @[control.py:95:Control.fir@130.4]
  assign _T_143 = _T_74 ? 3'h4 : _T_142; // @[control.py:95:Control.fir@131.4]
  assign _T_144 = _T_72 ? 3'h3 : _T_143; // @[control.py:95:Control.fir@132.4]
  assign _T_145 = _T_70 ? 3'h3 : _T_144; // @[control.py:95:Control.fir@133.4]
  assign _T_146 = _T_68 ? 3'h3 : _T_145; // @[control.py:95:Control.fir@134.4]
  assign _T_147 = _T_66 ? 3'h2 : _T_146; // @[control.py:95:Control.fir@135.4]
  assign _T_148 = _T_64 ? 3'h2 : _T_147; // @[control.py:95:Control.fir@136.4]
  assign _T_149 = _T_62 ? 3'h2 : _T_148; // @[control.py:95:Control.fir@137.4]
  assign _T_150 = _T_60 ? 3'h2 : _T_149; // @[control.py:95:Control.fir@138.4]
  assign _T_151 = _T_58 ? 3'h2 : _T_150; // @[control.py:95:Control.fir@139.4]
  assign _T_152 = _T_56 ? 3'h2 : _T_151; // @[control.py:95:Control.fir@140.4]
  assign _T_153 = _T_54 ? 3'h2 : _T_152; // @[control.py:95:Control.fir@141.4]
  assign _T_154 = _T_52 ? 3'h1 : _T_153; // @[control.py:95:Control.fir@142.4]
  assign _T_155 = _T_50 ? 3'h1 : _T_154; // @[control.py:95:Control.fir@143.4]
  assign _T_156 = _T_48 ? 3'h2 : _T_155; // @[control.py:95:Control.fir@144.4]
  assign _T_157 = _T_46 ? 3'h2 : _T_156; // @[control.py:95:Control.fir@145.4]
  assign _T_158 = _T_44 ? 3'h2 : _T_157; // @[control.py:95:Control.fir@146.4]
  assign _T_159 = _T_42 ? 3'h1 : _T_158; // @[control.py:95:Control.fir@147.4]
  assign _T_160 = _T_40 ? 3'h1 : _T_159; // @[control.py:95:Control.fir@148.4]
  assign _T_161 = _T_38 ? 3'h1 : _T_160; // @[control.py:95:Control.fir@149.4]
  assign _T_162 = _T_36 ? 3'h2 : _T_161; // @[control.py:95:Control.fir@150.4]
  assign _T_163 = _T_34 ? 3'h2 : _T_162; // @[control.py:95:Control.fir@151.4]
  assign _T_164 = _T_32 ? 3'h2 : _T_163; // @[control.py:95:Control.fir@152.4]
  assign _T_165 = _T_30 ? 3'h2 : _T_164; // @[control.py:95:Control.fir@153.4]
  assign _T_166 = _T_28 ? 3'h1 : _T_165; // @[control.py:95:Control.fir@154.4]
  assign _T_167 = _T_26 ? 3'h1 : _T_166; // @[control.py:95:Control.fir@155.4]
  assign _T_168 = _T_24 ? 3'h1 : _T_167; // @[control.py:95:Control.fir@156.4]
  assign _T_169 = _T_22 ? 3'h1 : _T_168; // @[control.py:95:Control.fir@157.4]
  assign _T_183 = _T_70 ? 1'h1 : _T_72; // @[control.py:95:Control.fir@171.4]
  assign _T_184 = _T_68 ? 1'h1 : _T_183; // @[control.py:95:Control.fir@172.4]
  assign _T_185 = _T_66 ? 1'h1 : _T_184; // @[control.py:95:Control.fir@173.4]
  assign _T_186 = _T_64 ? 1'h1 : _T_185; // @[control.py:95:Control.fir@174.4]
  assign _T_187 = _T_62 ? 1'h1 : _T_186; // @[control.py:95:Control.fir@175.4]
  assign _T_188 = _T_60 ? 1'h1 : _T_187; // @[control.py:95:Control.fir@176.4]
  assign _T_189 = _T_58 ? 1'h1 : _T_188; // @[control.py:95:Control.fir@177.4]
  assign _T_190 = _T_56 ? 1'h1 : _T_189; // @[control.py:95:Control.fir@178.4]
  assign _T_191 = _T_54 ? 1'h1 : _T_190; // @[control.py:95:Control.fir@179.4]
  assign _T_192 = _T_52 ? 1'h0 : _T_191; // @[control.py:95:Control.fir@180.4]
  assign _T_193 = _T_50 ? 1'h0 : _T_192; // @[control.py:95:Control.fir@181.4]
  assign _T_194 = _T_48 ? 1'h1 : _T_193; // @[control.py:95:Control.fir@182.4]
  assign _T_195 = _T_46 ? 1'h1 : _T_194; // @[control.py:95:Control.fir@183.4]
  assign _T_196 = _T_44 ? 1'h1 : _T_195; // @[control.py:95:Control.fir@184.4]
  assign _T_197 = _T_42 ? 1'h0 : _T_196; // @[control.py:95:Control.fir@185.4]
  assign _T_198 = _T_40 ? 1'h0 : _T_197; // @[control.py:95:Control.fir@186.4]
  assign _T_199 = _T_38 ? 1'h0 : _T_198; // @[control.py:95:Control.fir@187.4]
  assign _T_200 = _T_36 ? 1'h1 : _T_199; // @[control.py:95:Control.fir@188.4]
  assign _T_201 = _T_34 ? 1'h1 : _T_200; // @[control.py:95:Control.fir@189.4]
  assign _T_202 = _T_32 ? 1'h1 : _T_201; // @[control.py:95:Control.fir@190.4]
  assign _T_203 = _T_30 ? 1'h1 : _T_202; // @[control.py:95:Control.fir@191.4]
  assign _T_204 = _T_28 ? 1'h0 : _T_203; // @[control.py:95:Control.fir@192.4]
  assign _T_205 = _T_26 ? 1'h0 : _T_204; // @[control.py:95:Control.fir@193.4]
  assign _T_206 = _T_24 ? 1'h0 : _T_205; // @[control.py:95:Control.fir@194.4]
  assign _T_207 = _T_22 ? 1'h0 : _T_206; // @[control.py:95:Control.fir@195.4]
  assign _T_210 = _T_92 ? 5'h0 : 5'h10; // @[control.py:95:Control.fir@198.4]
  assign _T_211 = _T_90 ? 5'h0 : _T_210; // @[control.py:95:Control.fir@199.4]
  assign _T_212 = _T_88 ? 5'h0 : _T_211; // @[control.py:95:Control.fir@200.4]
  assign _T_213 = _T_86 ? 5'h0 : _T_212; // @[control.py:95:Control.fir@201.4]
  assign _T_214 = _T_84 ? 5'hf : _T_213; // @[control.py:95:Control.fir@202.4]
  assign _T_215 = _T_82 ? 5'he : _T_214; // @[control.py:95:Control.fir@203.4]
  assign _T_216 = _T_80 ? 5'hd : _T_215; // @[control.py:95:Control.fir@204.4]
  assign _T_217 = _T_78 ? 5'hc : _T_216; // @[control.py:95:Control.fir@205.4]
  assign _T_218 = _T_76 ? 5'hb : _T_217; // @[control.py:95:Control.fir@206.4]
  assign _T_219 = _T_74 ? 5'ha : _T_218; // @[control.py:95:Control.fir@207.4]
  assign _T_220 = _T_72 ? 5'h0 : _T_219; // @[control.py:95:Control.fir@208.4]
  assign _T_221 = _T_70 ? 5'h0 : _T_220; // @[control.py:95:Control.fir@209.4]
  assign _T_222 = _T_68 ? 5'h0 : _T_221; // @[control.py:95:Control.fir@210.4]
  assign _T_223 = _T_66 ? 5'h0 : _T_222; // @[control.py:95:Control.fir@211.4]
  assign _T_224 = _T_64 ? 5'h0 : _T_223; // @[control.py:95:Control.fir@212.4]
  assign _T_225 = _T_62 ? 5'h0 : _T_224; // @[control.py:95:Control.fir@213.4]
  assign _T_226 = _T_60 ? 5'h0 : _T_225; // @[control.py:95:Control.fir@214.4]
  assign _T_227 = _T_58 ? 5'h0 : _T_226; // @[control.py:95:Control.fir@215.4]
  assign _T_228 = _T_56 ? 5'h9 : _T_227; // @[control.py:95:Control.fir@216.4]
  assign _T_229 = _T_54 ? 5'h8 : _T_228; // @[control.py:95:Control.fir@217.4]
  assign _T_230 = _T_52 ? 5'h9 : _T_229; // @[control.py:95:Control.fir@218.4]
  assign _T_231 = _T_50 ? 5'h8 : _T_230; // @[control.py:95:Control.fir@219.4]
  assign _T_232 = _T_48 ? 5'h7 : _T_231; // @[control.py:95:Control.fir@220.4]
  assign _T_233 = _T_46 ? 5'h6 : _T_232; // @[control.py:95:Control.fir@221.4]
  assign _T_234 = _T_44 ? 5'h5 : _T_233; // @[control.py:95:Control.fir@222.4]
  assign _T_235 = _T_42 ? 5'h7 : _T_234; // @[control.py:95:Control.fir@223.4]
  assign _T_236 = _T_40 ? 5'h6 : _T_235; // @[control.py:95:Control.fir@224.4]
  assign _T_237 = _T_38 ? 5'h5 : _T_236; // @[control.py:95:Control.fir@225.4]
  assign _T_238 = _T_36 ? 5'h4 : _T_237; // @[control.py:95:Control.fir@226.4]
  assign _T_239 = _T_34 ? 5'h3 : _T_238; // @[control.py:95:Control.fir@227.4]
  assign _T_240 = _T_32 ? 5'h2 : _T_239; // @[control.py:95:Control.fir@228.4]
  assign _T_241 = _T_30 ? 5'h0 : _T_240; // @[control.py:95:Control.fir@229.4]
  assign _T_242 = _T_28 ? 5'h4 : _T_241; // @[control.py:95:Control.fir@230.4]
  assign _T_243 = _T_26 ? 5'h3 : _T_242; // @[control.py:95:Control.fir@231.4]
  assign _T_244 = _T_24 ? 5'h2 : _T_243; // @[control.py:95:Control.fir@232.4]
  assign _T_245 = _T_22 ? 5'h1 : _T_244; // @[control.py:95:Control.fir@233.4]
  assign _T_251 = _T_86 ? 1'h1 : _T_88; // @[control.py:95:Control.fir@239.4]
  assign _T_252 = _T_84 ? 1'h1 : _T_251; // @[control.py:95:Control.fir@240.4]
  assign _T_253 = _T_82 ? 1'h1 : _T_252; // @[control.py:95:Control.fir@241.4]
  assign _T_254 = _T_80 ? 1'h1 : _T_253; // @[control.py:95:Control.fir@242.4]
  assign _T_255 = _T_78 ? 1'h1 : _T_254; // @[control.py:95:Control.fir@243.4]
  assign _T_256 = _T_76 ? 1'h1 : _T_255; // @[control.py:95:Control.fir@244.4]
  assign _T_257 = _T_74 ? 1'h1 : _T_256; // @[control.py:95:Control.fir@245.4]
  assign _T_258 = _T_72 ? 1'h0 : _T_257; // @[control.py:95:Control.fir@246.4]
  assign _T_259 = _T_70 ? 1'h0 : _T_258; // @[control.py:95:Control.fir@247.4]
  assign _T_260 = _T_68 ? 1'h0 : _T_259; // @[control.py:95:Control.fir@248.4]
  assign _T_261 = _T_66 ? 1'h0 : _T_260; // @[control.py:95:Control.fir@249.4]
  assign _T_262 = _T_64 ? 1'h0 : _T_261; // @[control.py:95:Control.fir@250.4]
  assign _T_263 = _T_62 ? 1'h0 : _T_262; // @[control.py:95:Control.fir@251.4]
  assign _T_264 = _T_60 ? 1'h0 : _T_263; // @[control.py:95:Control.fir@252.4]
  assign _T_265 = _T_58 ? 1'h0 : _T_264; // @[control.py:95:Control.fir@253.4]
  assign _T_266 = _T_56 ? 1'h0 : _T_265; // @[control.py:95:Control.fir@254.4]
  assign _T_267 = _T_54 ? 1'h0 : _T_266; // @[control.py:95:Control.fir@255.4]
  assign _T_268 = _T_52 ? 1'h0 : _T_267; // @[control.py:95:Control.fir@256.4]
  assign _T_269 = _T_50 ? 1'h0 : _T_268; // @[control.py:95:Control.fir@257.4]
  assign _T_270 = _T_48 ? 1'h0 : _T_269; // @[control.py:95:Control.fir@258.4]
  assign _T_271 = _T_46 ? 1'h0 : _T_270; // @[control.py:95:Control.fir@259.4]
  assign _T_272 = _T_44 ? 1'h0 : _T_271; // @[control.py:95:Control.fir@260.4]
  assign _T_273 = _T_42 ? 1'h0 : _T_272; // @[control.py:95:Control.fir@261.4]
  assign _T_274 = _T_40 ? 1'h0 : _T_273; // @[control.py:95:Control.fir@262.4]
  assign _T_275 = _T_38 ? 1'h0 : _T_274; // @[control.py:95:Control.fir@263.4]
  assign _T_276 = _T_36 ? 1'h0 : _T_275; // @[control.py:95:Control.fir@264.4]
  assign _T_277 = _T_34 ? 1'h0 : _T_276; // @[control.py:95:Control.fir@265.4]
  assign _T_278 = _T_32 ? 1'h0 : _T_277; // @[control.py:95:Control.fir@266.4]
  assign _T_279 = _T_30 ? 1'h0 : _T_278; // @[control.py:95:Control.fir@267.4]
  assign _T_280 = _T_28 ? 1'h0 : _T_279; // @[control.py:95:Control.fir@268.4]
  assign _T_281 = _T_26 ? 1'h0 : _T_280; // @[control.py:95:Control.fir@269.4]
  assign _T_282 = _T_24 ? 1'h0 : _T_281; // @[control.py:95:Control.fir@270.4]
  assign _T_283 = _T_22 ? 1'h0 : _T_282; // @[control.py:95:Control.fir@271.4]
  assign _T_289 = _T_86 ? 1'h0 : _T_88; // @[control.py:95:Control.fir@277.4]
  assign _T_290 = _T_84 ? 1'h0 : _T_289; // @[control.py:95:Control.fir@278.4]
  assign _T_291 = _T_82 ? 1'h0 : _T_290; // @[control.py:95:Control.fir@279.4]
  assign _T_292 = _T_80 ? 1'h0 : _T_291; // @[control.py:95:Control.fir@280.4]
  assign _T_293 = _T_78 ? 1'h0 : _T_292; // @[control.py:95:Control.fir@281.4]
  assign _T_294 = _T_76 ? 1'h0 : _T_293; // @[control.py:95:Control.fir@282.4]
  assign _T_295 = _T_74 ? 1'h0 : _T_294; // @[control.py:95:Control.fir@283.4]
  assign _T_296 = _T_72 ? 1'h0 : _T_295; // @[control.py:95:Control.fir@284.4]
  assign _T_297 = _T_70 ? 1'h0 : _T_296; // @[control.py:95:Control.fir@285.4]
  assign _T_298 = _T_68 ? 1'h0 : _T_297; // @[control.py:95:Control.fir@286.4]
  assign _T_299 = _T_66 ? 1'h0 : _T_298; // @[control.py:95:Control.fir@287.4]
  assign _T_300 = _T_64 ? 1'h0 : _T_299; // @[control.py:95:Control.fir@288.4]
  assign _T_301 = _T_62 ? 1'h0 : _T_300; // @[control.py:95:Control.fir@289.4]
  assign _T_302 = _T_60 ? 1'h0 : _T_301; // @[control.py:95:Control.fir@290.4]
  assign _T_303 = _T_58 ? 1'h0 : _T_302; // @[control.py:95:Control.fir@291.4]
  assign _T_304 = _T_56 ? 1'h0 : _T_303; // @[control.py:95:Control.fir@292.4]
  assign _T_305 = _T_54 ? 1'h0 : _T_304; // @[control.py:95:Control.fir@293.4]
  assign _T_306 = _T_52 ? 1'h0 : _T_305; // @[control.py:95:Control.fir@294.4]
  assign _T_307 = _T_50 ? 1'h0 : _T_306; // @[control.py:95:Control.fir@295.4]
  assign _T_308 = _T_48 ? 1'h0 : _T_307; // @[control.py:95:Control.fir@296.4]
  assign _T_309 = _T_46 ? 1'h0 : _T_308; // @[control.py:95:Control.fir@297.4]
  assign _T_310 = _T_44 ? 1'h0 : _T_309; // @[control.py:95:Control.fir@298.4]
  assign _T_311 = _T_42 ? 1'h0 : _T_310; // @[control.py:95:Control.fir@299.4]
  assign _T_312 = _T_40 ? 1'h0 : _T_311; // @[control.py:95:Control.fir@300.4]
  assign _T_313 = _T_38 ? 1'h0 : _T_312; // @[control.py:95:Control.fir@301.4]
  assign _T_314 = _T_36 ? 1'h0 : _T_313; // @[control.py:95:Control.fir@302.4]
  assign _T_315 = _T_34 ? 1'h0 : _T_314; // @[control.py:95:Control.fir@303.4]
  assign _T_316 = _T_32 ? 1'h0 : _T_315; // @[control.py:95:Control.fir@304.4]
  assign _T_317 = _T_30 ? 1'h0 : _T_316; // @[control.py:95:Control.fir@305.4]
  assign _T_318 = _T_28 ? 1'h0 : _T_317; // @[control.py:95:Control.fir@306.4]
  assign _T_319 = _T_26 ? 1'h0 : _T_318; // @[control.py:95:Control.fir@307.4]
  assign _T_320 = _T_24 ? 1'h0 : _T_319; // @[control.py:95:Control.fir@308.4]
  assign _T_321 = _T_22 ? 1'h0 : _T_320; // @[control.py:95:Control.fir@309.4]
  assign _T_338 = _T_64 ? 1'h1 : _T_66; // @[control.py:95:Control.fir@326.4]
  assign _T_339 = _T_62 ? 1'h1 : _T_338; // @[control.py:95:Control.fir@327.4]
  assign _T_340 = _T_60 ? 1'h1 : _T_339; // @[control.py:95:Control.fir@328.4]
  assign _T_341 = _T_58 ? 1'h1 : _T_340; // @[control.py:95:Control.fir@329.4]
  assign _T_342 = _T_56 ? 1'h0 : _T_341; // @[control.py:95:Control.fir@330.4]
  assign _T_343 = _T_54 ? 1'h0 : _T_342; // @[control.py:95:Control.fir@331.4]
  assign _T_344 = _T_52 ? 1'h0 : _T_343; // @[control.py:95:Control.fir@332.4]
  assign _T_345 = _T_50 ? 1'h0 : _T_344; // @[control.py:95:Control.fir@333.4]
  assign _T_346 = _T_48 ? 1'h0 : _T_345; // @[control.py:95:Control.fir@334.4]
  assign _T_347 = _T_46 ? 1'h0 : _T_346; // @[control.py:95:Control.fir@335.4]
  assign _T_348 = _T_44 ? 1'h0 : _T_347; // @[control.py:95:Control.fir@336.4]
  assign _T_349 = _T_42 ? 1'h0 : _T_348; // @[control.py:95:Control.fir@337.4]
  assign _T_350 = _T_40 ? 1'h0 : _T_349; // @[control.py:95:Control.fir@338.4]
  assign _T_351 = _T_38 ? 1'h0 : _T_350; // @[control.py:95:Control.fir@339.4]
  assign _T_352 = _T_36 ? 1'h0 : _T_351; // @[control.py:95:Control.fir@340.4]
  assign _T_353 = _T_34 ? 1'h0 : _T_352; // @[control.py:95:Control.fir@341.4]
  assign _T_354 = _T_32 ? 1'h0 : _T_353; // @[control.py:95:Control.fir@342.4]
  assign _T_355 = _T_30 ? 1'h0 : _T_354; // @[control.py:95:Control.fir@343.4]
  assign _T_356 = _T_28 ? 1'h0 : _T_355; // @[control.py:95:Control.fir@344.4]
  assign _T_357 = _T_26 ? 1'h0 : _T_356; // @[control.py:95:Control.fir@345.4]
  assign _T_358 = _T_24 ? 1'h0 : _T_357; // @[control.py:95:Control.fir@346.4]
  assign _T_359 = _T_22 ? 1'h0 : _T_358; // @[control.py:95:Control.fir@347.4]
  assign _T_375 = _T_66 ? 1'h0 : _T_184; // @[control.py:95:Control.fir@363.4]
  assign _T_376 = _T_64 ? 1'h0 : _T_375; // @[control.py:95:Control.fir@364.4]
  assign _T_377 = _T_62 ? 1'h0 : _T_376; // @[control.py:95:Control.fir@365.4]
  assign _T_378 = _T_60 ? 1'h0 : _T_377; // @[control.py:95:Control.fir@366.4]
  assign _T_379 = _T_58 ? 1'h0 : _T_378; // @[control.py:95:Control.fir@367.4]
  assign _T_380 = _T_56 ? 1'h0 : _T_379; // @[control.py:95:Control.fir@368.4]
  assign _T_381 = _T_54 ? 1'h0 : _T_380; // @[control.py:95:Control.fir@369.4]
  assign _T_382 = _T_52 ? 1'h0 : _T_381; // @[control.py:95:Control.fir@370.4]
  assign _T_383 = _T_50 ? 1'h0 : _T_382; // @[control.py:95:Control.fir@371.4]
  assign _T_384 = _T_48 ? 1'h0 : _T_383; // @[control.py:95:Control.fir@372.4]
  assign _T_385 = _T_46 ? 1'h0 : _T_384; // @[control.py:95:Control.fir@373.4]
  assign _T_386 = _T_44 ? 1'h0 : _T_385; // @[control.py:95:Control.fir@374.4]
  assign _T_387 = _T_42 ? 1'h0 : _T_386; // @[control.py:95:Control.fir@375.4]
  assign _T_388 = _T_40 ? 1'h0 : _T_387; // @[control.py:95:Control.fir@376.4]
  assign _T_389 = _T_38 ? 1'h0 : _T_388; // @[control.py:95:Control.fir@377.4]
  assign _T_390 = _T_36 ? 1'h0 : _T_389; // @[control.py:95:Control.fir@378.4]
  assign _T_391 = _T_34 ? 1'h0 : _T_390; // @[control.py:95:Control.fir@379.4]
  assign _T_392 = _T_32 ? 1'h0 : _T_391; // @[control.py:95:Control.fir@380.4]
  assign _T_393 = _T_30 ? 1'h0 : _T_392; // @[control.py:95:Control.fir@381.4]
  assign _T_394 = _T_28 ? 1'h0 : _T_393; // @[control.py:95:Control.fir@382.4]
  assign _T_395 = _T_26 ? 1'h0 : _T_394; // @[control.py:95:Control.fir@383.4]
  assign _T_396 = _T_24 ? 1'h0 : _T_395; // @[control.py:95:Control.fir@384.4]
  assign _T_397 = _T_22 ? 1'h0 : _T_396; // @[control.py:95:Control.fir@385.4]
  assign _T_410 = _T_72 ? 2'h2 : 2'h0; // @[control.py:95:Control.fir@398.4]
  assign _T_411 = _T_70 ? 2'h1 : _T_410; // @[control.py:95:Control.fir@399.4]
  assign _T_412 = _T_68 ? 2'h0 : _T_411; // @[control.py:95:Control.fir@400.4]
  assign _T_413 = _T_66 ? 2'h2 : _T_412; // @[control.py:95:Control.fir@401.4]
  assign _T_414 = _T_64 ? 2'h1 : _T_413; // @[control.py:95:Control.fir@402.4]
  assign _T_415 = _T_62 ? 2'h2 : _T_414; // @[control.py:95:Control.fir@403.4]
  assign _T_416 = _T_60 ? 2'h1 : _T_415; // @[control.py:95:Control.fir@404.4]
  assign _T_417 = _T_58 ? 2'h0 : _T_416; // @[control.py:95:Control.fir@405.4]
  assign _T_418 = _T_56 ? 2'h0 : _T_417; // @[control.py:95:Control.fir@406.4]
  assign _T_419 = _T_54 ? 2'h0 : _T_418; // @[control.py:95:Control.fir@407.4]
  assign _T_420 = _T_52 ? 2'h0 : _T_419; // @[control.py:95:Control.fir@408.4]
  assign _T_421 = _T_50 ? 2'h0 : _T_420; // @[control.py:95:Control.fir@409.4]
  assign _T_422 = _T_48 ? 2'h0 : _T_421; // @[control.py:95:Control.fir@410.4]
  assign _T_423 = _T_46 ? 2'h0 : _T_422; // @[control.py:95:Control.fir@411.4]
  assign _T_424 = _T_44 ? 2'h0 : _T_423; // @[control.py:95:Control.fir@412.4]
  assign _T_425 = _T_42 ? 2'h0 : _T_424; // @[control.py:95:Control.fir@413.4]
  assign _T_426 = _T_40 ? 2'h0 : _T_425; // @[control.py:95:Control.fir@414.4]
  assign _T_427 = _T_38 ? 2'h0 : _T_426; // @[control.py:95:Control.fir@415.4]
  assign _T_428 = _T_36 ? 2'h0 : _T_427; // @[control.py:95:Control.fir@416.4]
  assign _T_429 = _T_34 ? 2'h0 : _T_428; // @[control.py:95:Control.fir@417.4]
  assign _T_430 = _T_32 ? 2'h0 : _T_429; // @[control.py:95:Control.fir@418.4]
  assign _T_431 = _T_30 ? 2'h0 : _T_430; // @[control.py:95:Control.fir@419.4]
  assign _T_432 = _T_28 ? 2'h0 : _T_431; // @[control.py:95:Control.fir@420.4]
  assign _T_433 = _T_26 ? 2'h0 : _T_432; // @[control.py:95:Control.fir@421.4]
  assign _T_434 = _T_24 ? 2'h0 : _T_433; // @[control.py:95:Control.fir@422.4]
  assign _T_435 = _T_22 ? 2'h0 : _T_434; // @[control.py:95:Control.fir@423.4]
  assign _T_453 = _T_62 ? 1'h0 : _T_338; // @[control.py:95:Control.fir@441.4]
  assign _T_454 = _T_60 ? 1'h0 : _T_453; // @[control.py:95:Control.fir@442.4]
  assign _T_455 = _T_58 ? 1'h0 : _T_454; // @[control.py:95:Control.fir@443.4]
  assign _T_456 = _T_56 ? 1'h0 : _T_455; // @[control.py:95:Control.fir@444.4]
  assign _T_457 = _T_54 ? 1'h0 : _T_456; // @[control.py:95:Control.fir@445.4]
  assign _T_458 = _T_52 ? 1'h0 : _T_457; // @[control.py:95:Control.fir@446.4]
  assign _T_459 = _T_50 ? 1'h0 : _T_458; // @[control.py:95:Control.fir@447.4]
  assign _T_460 = _T_48 ? 1'h0 : _T_459; // @[control.py:95:Control.fir@448.4]
  assign _T_461 = _T_46 ? 1'h0 : _T_460; // @[control.py:95:Control.fir@449.4]
  assign _T_462 = _T_44 ? 1'h0 : _T_461; // @[control.py:95:Control.fir@450.4]
  assign _T_463 = _T_42 ? 1'h0 : _T_462; // @[control.py:95:Control.fir@451.4]
  assign _T_464 = _T_40 ? 1'h0 : _T_463; // @[control.py:95:Control.fir@452.4]
  assign _T_465 = _T_38 ? 1'h0 : _T_464; // @[control.py:95:Control.fir@453.4]
  assign _T_466 = _T_36 ? 1'h0 : _T_465; // @[control.py:95:Control.fir@454.4]
  assign _T_467 = _T_34 ? 1'h0 : _T_466; // @[control.py:95:Control.fir@455.4]
  assign _T_468 = _T_32 ? 1'h0 : _T_467; // @[control.py:95:Control.fir@456.4]
  assign _T_469 = _T_30 ? 1'h0 : _T_468; // @[control.py:95:Control.fir@457.4]
  assign _T_470 = _T_28 ? 1'h0 : _T_469; // @[control.py:95:Control.fir@458.4]
  assign _T_471 = _T_26 ? 1'h0 : _T_470; // @[control.py:95:Control.fir@459.4]
  assign _T_472 = _T_24 ? 1'h0 : _T_471; // @[control.py:95:Control.fir@460.4]
  assign _T_473 = _T_22 ? 1'h0 : _T_472; // @[control.py:95:Control.fir@461.4]
  assign _T_476 = _T_92 ? 3'h4 : 3'h0; // @[control.py:95:Control.fir@464.4]
  assign _T_477 = _T_90 ? 3'h3 : _T_476; // @[control.py:95:Control.fir@465.4]
  assign _T_478 = _T_88 ? 3'h2 : _T_477; // @[control.py:95:Control.fir@466.4]
  assign _T_479 = _T_86 ? 3'h2 : _T_478; // @[control.py:95:Control.fir@467.4]
  assign _T_480 = _T_84 ? 3'h0 : _T_479; // @[control.py:95:Control.fir@468.4]
  assign _T_481 = _T_82 ? 3'h0 : _T_480; // @[control.py:95:Control.fir@469.4]
  assign _T_482 = _T_80 ? 3'h0 : _T_481; // @[control.py:95:Control.fir@470.4]
  assign _T_483 = _T_78 ? 3'h0 : _T_482; // @[control.py:95:Control.fir@471.4]
  assign _T_484 = _T_76 ? 3'h0 : _T_483; // @[control.py:95:Control.fir@472.4]
  assign _T_485 = _T_74 ? 3'h0 : _T_484; // @[control.py:95:Control.fir@473.4]
  assign _T_486 = _T_72 ? 3'h0 : _T_485; // @[control.py:95:Control.fir@474.4]
  assign _T_487 = _T_70 ? 3'h0 : _T_486; // @[control.py:95:Control.fir@475.4]
  assign _T_488 = _T_68 ? 3'h0 : _T_487; // @[control.py:95:Control.fir@476.4]
  assign _T_489 = _T_66 ? 3'h1 : _T_488; // @[control.py:95:Control.fir@477.4]
  assign _T_490 = _T_64 ? 3'h1 : _T_489; // @[control.py:95:Control.fir@478.4]
  assign _T_491 = _T_62 ? 3'h1 : _T_490; // @[control.py:95:Control.fir@479.4]
  assign _T_492 = _T_60 ? 3'h1 : _T_491; // @[control.py:95:Control.fir@480.4]
  assign _T_493 = _T_58 ? 3'h1 : _T_492; // @[control.py:95:Control.fir@481.4]
  assign _T_494 = _T_56 ? 3'h0 : _T_493; // @[control.py:95:Control.fir@482.4]
  assign _T_495 = _T_54 ? 3'h0 : _T_494; // @[control.py:95:Control.fir@483.4]
  assign _T_496 = _T_52 ? 3'h0 : _T_495; // @[control.py:95:Control.fir@484.4]
  assign _T_497 = _T_50 ? 3'h0 : _T_496; // @[control.py:95:Control.fir@485.4]
  assign _T_498 = _T_48 ? 3'h0 : _T_497; // @[control.py:95:Control.fir@486.4]
  assign _T_499 = _T_46 ? 3'h0 : _T_498; // @[control.py:95:Control.fir@487.4]
  assign _T_500 = _T_44 ? 3'h0 : _T_499; // @[control.py:95:Control.fir@488.4]
  assign _T_501 = _T_42 ? 3'h0 : _T_500; // @[control.py:95:Control.fir@489.4]
  assign _T_502 = _T_40 ? 3'h0 : _T_501; // @[control.py:95:Control.fir@490.4]
  assign _T_503 = _T_38 ? 3'h0 : _T_502; // @[control.py:95:Control.fir@491.4]
  assign _T_504 = _T_36 ? 3'h0 : _T_503; // @[control.py:95:Control.fir@492.4]
  assign _T_505 = _T_34 ? 3'h0 : _T_504; // @[control.py:95:Control.fir@493.4]
  assign _T_506 = _T_32 ? 3'h0 : _T_505; // @[control.py:95:Control.fir@494.4]
  assign _T_507 = _T_30 ? 3'h0 : _T_506; // @[control.py:95:Control.fir@495.4]
  assign _T_508 = _T_28 ? 3'h0 : _T_507; // @[control.py:95:Control.fir@496.4]
  assign _T_509 = _T_26 ? 3'h0 : _T_508; // @[control.py:95:Control.fir@497.4]
  assign _T_510 = _T_24 ? 3'h0 : _T_509; // @[control.py:95:Control.fir@498.4]
  assign _T_511 = _T_22 ? 3'h0 : _T_510; // @[control.py:95:Control.fir@499.4]
  assign _T_518 = _T_84 ? 1'h0 : _T_251; // @[control.py:95:Control.fir@506.4]
  assign _T_519 = _T_82 ? 1'h0 : _T_518; // @[control.py:95:Control.fir@507.4]
  assign _T_520 = _T_80 ? 1'h0 : _T_519; // @[control.py:95:Control.fir@508.4]
  assign _T_521 = _T_78 ? 1'h0 : _T_520; // @[control.py:95:Control.fir@509.4]
  assign _T_522 = _T_76 ? 1'h0 : _T_521; // @[control.py:95:Control.fir@510.4]
  assign _T_523 = _T_74 ? 1'h0 : _T_522; // @[control.py:95:Control.fir@511.4]
  assign _T_524 = _T_72 ? 1'h0 : _T_523; // @[control.py:95:Control.fir@512.4]
  assign _T_525 = _T_70 ? 1'h0 : _T_524; // @[control.py:95:Control.fir@513.4]
  assign _T_526 = _T_68 ? 1'h0 : _T_525; // @[control.py:95:Control.fir@514.4]
  assign _T_527 = _T_66 ? 1'h0 : _T_526; // @[control.py:95:Control.fir@515.4]
  assign _T_528 = _T_64 ? 1'h0 : _T_527; // @[control.py:95:Control.fir@516.4]
  assign _T_529 = _T_62 ? 1'h0 : _T_528; // @[control.py:95:Control.fir@517.4]
  assign _T_530 = _T_60 ? 1'h0 : _T_529; // @[control.py:95:Control.fir@518.4]
  assign _T_531 = _T_58 ? 1'h0 : _T_530; // @[control.py:95:Control.fir@519.4]
  assign _T_532 = _T_56 ? 1'h0 : _T_531; // @[control.py:95:Control.fir@520.4]
  assign _T_533 = _T_54 ? 1'h0 : _T_532; // @[control.py:95:Control.fir@521.4]
  assign _T_534 = _T_52 ? 1'h0 : _T_533; // @[control.py:95:Control.fir@522.4]
  assign _T_535 = _T_50 ? 1'h0 : _T_534; // @[control.py:95:Control.fir@523.4]
  assign _T_536 = _T_48 ? 1'h0 : _T_535; // @[control.py:95:Control.fir@524.4]
  assign _T_537 = _T_46 ? 1'h0 : _T_536; // @[control.py:95:Control.fir@525.4]
  assign _T_538 = _T_44 ? 1'h0 : _T_537; // @[control.py:95:Control.fir@526.4]
  assign _T_539 = _T_42 ? 1'h0 : _T_538; // @[control.py:95:Control.fir@527.4]
  assign _T_540 = _T_40 ? 1'h0 : _T_539; // @[control.py:95:Control.fir@528.4]
  assign _T_541 = _T_38 ? 1'h0 : _T_540; // @[control.py:95:Control.fir@529.4]
  assign _T_542 = _T_36 ? 1'h0 : _T_541; // @[control.py:95:Control.fir@530.4]
  assign _T_543 = _T_34 ? 1'h0 : _T_542; // @[control.py:95:Control.fir@531.4]
  assign _T_544 = _T_32 ? 1'h0 : _T_543; // @[control.py:95:Control.fir@532.4]
  assign _T_545 = _T_30 ? 1'h0 : _T_544; // @[control.py:95:Control.fir@533.4]
  assign _T_546 = _T_28 ? 1'h0 : _T_545; // @[control.py:95:Control.fir@534.4]
  assign _T_547 = _T_26 ? 1'h0 : _T_546; // @[control.py:95:Control.fir@535.4]
  assign _T_548 = _T_24 ? 1'h0 : _T_547; // @[control.py:95:Control.fir@536.4]
  assign _T_549 = _T_22 ? 1'h0 : _T_548; // @[control.py:95:Control.fir@537.4]
  assign io_ctrl_Reg_Write = _T_20 ? 1'h1 : _T_131; // @[control.py:114:Control.fir@549.4]
  assign io_ctrl_Imm_Sel = _T_20 ? 3'h1 : _T_169; // @[control.py:98:Control.fir@539.4]
  assign io_ctrl_ALU_Src = _T_20 ? 1'h0 : _T_207; // @[control.py:101:Control.fir@540.4]
  assign io_ctrl_ALUOp = _T_20 ? 5'h0 : _T_245; // @[control.py:102:Control.fir@541.4]
  assign io_ctrl_Branch = _T_20 ? 1'h0 : _T_283; // @[control.py:103:Control.fir@542.4]
  assign io_ctrl_Branch_Src = _T_20 ? 1'h0 : _T_321; // @[control.py:104:Control.fir@543.4]
  assign io_ctrl_Mem_Read = _T_20 ? 1'h0 : _T_359; // @[control.py:108:Control.fir@545.4]
  assign io_ctrl_Mem_Write = _T_20 ? 1'h0 : _T_397; // @[control.py:109:Control.fir@546.4]
  assign io_ctrl_Data_Size = _T_20 ? 2'h0 : _T_435; // @[control.py:110:Control.fir@547.4]
  assign io_ctrl_Load_Type = _T_20 ? 1'h0 : _T_473; // @[control.py:111:Control.fir@548.4]
  assign io_ctrl_Mem_to_Reg = _T_20 ? 3'h0 : _T_511; // @[control.py:115:Control.fir@550.4]
  assign io_ctrl_Jump_Type = _T_20 ? 1'h0 : _T_549; // @[control.py:105:Control.fir@544.4]
endmodule
