module ALU( // @[alu.py:21:ALU.fir@2.2]
  input         clock, // @[rawmodule.py:100:ALU.fir@3.4]
  input         reset, // @[rawmodule.py:101:ALU.fir@4.4]
  input  [31:0] io_src_a, // @[alu.py:11:ALU.fir@5.4]
  input  [31:0] io_src_b, // @[alu.py:11:ALU.fir@5.4]
  input  [4:0]  io_ALUOp, // @[alu.py:11:ALU.fir@5.4]
  output [31:0] io_sum, // @[alu.py:11:ALU.fir@5.4]
  output        io_conflag // @[alu.py:11:ALU.fir@5.4]
);
  wire [5:0] _T_9; // @[alu.py:24:ALU.fir@7.4]
  wire [32:0] _T_10; // @[alu.py:26:ALU.fir@8.4]
  wire [32:0] _T_11; // @[alu.py:27:ALU.fir@9.4]
  wire [31:0] _T_12; // @[alu.py:28:ALU.fir@10.4]
  wire [31:0] _T_13; // @[alu.py:29:ALU.fir@11.4]
  wire [31:0] _T_14; // @[alu.py:30:ALU.fir@12.4]
  wire [94:0] _GEN_0; // @[alu.py:31:ALU.fir@13.4]
  wire [94:0] _T_15; // @[alu.py:31:ALU.fir@13.4]
  wire [31:0] _T_16; // @[alu.py:32:ALU.fir@14.4]
  wire [31:0] _T_17; // @[alu.py:33:ALU.fir@15.4]
  wire [31:0] _T_18; // @[alu.py:33:ALU.fir@16.4]
  wire [31:0] _T_19; // @[alu.py:33:ALU.fir@17.4]
  wire [31:0] _T_21; // @[alu.py:34:ALU.fir@19.4]
  wire  _T_22; // @[alu.py:34:ALU.fir@20.4]
  wire  _T_23; // @[alu.py:35:ALU.fir@21.4]
  wire  _T_24; // @[mux.py:72:ALU.fir@22.4]
  wire [31:0] _T_25; // @[alu.py:35:ALU.fir@23.4]
  wire  _T_26; // @[mux.py:72:ALU.fir@24.4]
  wire [31:0] _T_27; // @[alu.py:35:ALU.fir@25.4]
  wire  _T_28; // @[mux.py:72:ALU.fir@26.4]
  wire [31:0] _T_29; // @[alu.py:35:ALU.fir@27.4]
  wire  _T_30; // @[mux.py:72:ALU.fir@28.4]
  wire [31:0] _T_31; // @[alu.py:35:ALU.fir@29.4]
  wire  _T_32; // @[mux.py:72:ALU.fir@30.4]
  wire [94:0] _T_33; // @[alu.py:35:ALU.fir@31.4]
  wire  _T_34; // @[mux.py:72:ALU.fir@32.4]
  wire [94:0] _T_35; // @[alu.py:35:ALU.fir@33.4]
  wire  _T_36; // @[mux.py:72:ALU.fir@34.4]
  wire [94:0] _T_37; // @[alu.py:35:ALU.fir@35.4]
  wire  _T_38; // @[mux.py:72:ALU.fir@36.4]
  wire [94:0] _T_39; // @[alu.py:35:ALU.fir@37.4]
  wire  _T_40; // @[mux.py:72:ALU.fir@38.4]
  wire [94:0] _T_41; // @[alu.py:35:ALU.fir@39.4]
  wire  _T_42; // @[mux.py:72:ALU.fir@40.4]
  wire [94:0] _T_43; // @[alu.py:35:ALU.fir@41.4]
  wire  _T_46; // @[alu.py:39:ALU.fir@45.4]
  wire  _T_55; // @[alu.py:42:ALU.fir@54.4]
  wire  _T_57; // @[alu.py:44:ALU.fir@56.4]
  wire  _T_58; // @[mux.py:72:ALU.fir@57.4]
  wire  _T_59; // @[alu.py:44:ALU.fir@58.4]
  wire  _T_60; // @[mux.py:72:ALU.fir@59.4]
  wire  _T_61; // @[alu.py:44:ALU.fir@60.4]
  wire  _T_62; // @[mux.py:72:ALU.fir@61.4]
  wire  _T_63; // @[alu.py:44:ALU.fir@62.4]
  wire  _T_64; // @[mux.py:72:ALU.fir@63.4]
  wire  _T_65; // @[alu.py:44:ALU.fir@64.4]
  wire  _T_66; // @[mux.py:72:ALU.fir@65.4]
  wire  _T_67; // @[alu.py:44:ALU.fir@66.4]
  wire  _T_68; // @[mux.py:72:ALU.fir@67.4]
  assign _T_9 = io_src_b[5:0]; // @[alu.py:24:ALU.fir@7.4]
  assign _T_10 = io_src_a + io_src_b; // @[alu.py:26:ALU.fir@8.4]
  assign _T_11 = io_src_a - io_src_b; // @[alu.py:27:ALU.fir@9.4]
  assign _T_12 = io_src_a & io_src_b; // @[alu.py:28:ALU.fir@10.4]
  assign _T_13 = io_src_a | io_src_b; // @[alu.py:29:ALU.fir@11.4]
  assign _T_14 = io_src_a ^ io_src_b; // @[alu.py:30:ALU.fir@12.4]
  assign _GEN_0 = {{63'd0}, io_src_a}; // @[alu.py:31:ALU.fir@13.4]
  assign _T_15 = _GEN_0 << _T_9; // @[alu.py:31:ALU.fir@13.4]
  assign _T_16 = io_src_a >> _T_9; // @[alu.py:32:ALU.fir@14.4]
  assign _T_17 = $signed(io_src_a); // @[alu.py:33:ALU.fir@15.4]
  assign _T_18 = $signed(_T_17) >>> _T_9; // @[alu.py:33:ALU.fir@16.4]
  assign _T_19 = $unsigned(_T_18); // @[alu.py:33:ALU.fir@17.4]
  assign _T_21 = $signed(io_src_b); // @[alu.py:34:ALU.fir@19.4]
  assign _T_22 = $signed(_T_17) < $signed(_T_21); // @[alu.py:34:ALU.fir@20.4]
  assign _T_23 = io_src_a < io_src_b; // @[alu.py:35:ALU.fir@21.4]
  assign _T_24 = io_ALUOp == 5'h9; // @[mux.py:72:ALU.fir@22.4]
  assign _T_25 = _T_24 ? {{31'd0}, _T_23} : io_src_b; // @[alu.py:35:ALU.fir@23.4]
  assign _T_26 = io_ALUOp == 5'h8; // @[mux.py:72:ALU.fir@24.4]
  assign _T_27 = _T_26 ? {{31'd0}, _T_22} : _T_25; // @[alu.py:35:ALU.fir@25.4]
  assign _T_28 = io_ALUOp == 5'h7; // @[mux.py:72:ALU.fir@26.4]
  assign _T_29 = _T_28 ? _T_19 : _T_27; // @[alu.py:35:ALU.fir@27.4]
  assign _T_30 = io_ALUOp == 5'h6; // @[mux.py:72:ALU.fir@28.4]
  assign _T_31 = _T_30 ? _T_16 : _T_29; // @[alu.py:35:ALU.fir@29.4]
  assign _T_32 = io_ALUOp == 5'h5; // @[mux.py:72:ALU.fir@30.4]
  assign _T_33 = _T_32 ? _T_15 : {{63'd0}, _T_31}; // @[alu.py:35:ALU.fir@31.4]
  assign _T_34 = io_ALUOp == 5'h4; // @[mux.py:72:ALU.fir@32.4]
  assign _T_35 = _T_34 ? {{63'd0}, _T_14} : _T_33; // @[alu.py:35:ALU.fir@33.4]
  assign _T_36 = io_ALUOp == 5'h3; // @[mux.py:72:ALU.fir@34.4]
  assign _T_37 = _T_36 ? {{63'd0}, _T_13} : _T_35; // @[alu.py:35:ALU.fir@35.4]
  assign _T_38 = io_ALUOp == 5'h2; // @[mux.py:72:ALU.fir@36.4]
  assign _T_39 = _T_38 ? {{63'd0}, _T_12} : _T_37; // @[alu.py:35:ALU.fir@37.4]
  assign _T_40 = io_ALUOp == 5'h1; // @[mux.py:72:ALU.fir@38.4]
  assign _T_41 = _T_40 ? {{62'd0}, _T_11} : _T_39; // @[alu.py:35:ALU.fir@39.4]
  assign _T_42 = io_ALUOp == 5'h0; // @[mux.py:72:ALU.fir@40.4]
  assign _T_43 = _T_42 ? {{62'd0}, _T_10} : _T_41; // @[alu.py:35:ALU.fir@41.4]
  assign _T_46 = $signed(_T_17) == $signed(_T_21); // @[alu.py:39:ALU.fir@45.4]
  assign _T_55 = $signed(_T_17) >= $signed(_T_21); // @[alu.py:42:ALU.fir@54.4]
  assign _T_57 = io_src_a >= io_src_b; // @[alu.py:44:ALU.fir@56.4]
  assign _T_58 = io_ALUOp == 5'hf; // @[mux.py:72:ALU.fir@57.4]
  assign _T_59 = _T_58 ? _T_57 : 1'h0; // @[alu.py:44:ALU.fir@58.4]
  assign _T_60 = io_ALUOp == 5'he; // @[mux.py:72:ALU.fir@59.4]
  assign _T_61 = _T_60 ? _T_23 : _T_59; // @[alu.py:44:ALU.fir@60.4]
  assign _T_62 = io_ALUOp == 5'hd; // @[mux.py:72:ALU.fir@61.4]
  assign _T_63 = _T_62 ? _T_55 : _T_61; // @[alu.py:44:ALU.fir@62.4]
  assign _T_64 = io_ALUOp == 5'hc; // @[mux.py:72:ALU.fir@63.4]
  assign _T_65 = _T_64 ? _T_22 : _T_63; // @[alu.py:44:ALU.fir@64.4]
  assign _T_66 = io_ALUOp == 5'hb; // @[mux.py:72:ALU.fir@65.4]
  assign _T_67 = _T_66 ? _T_46 : _T_65; // @[alu.py:44:ALU.fir@66.4]
  assign _T_68 = io_ALUOp == 5'ha; // @[mux.py:72:ALU.fir@67.4]
  assign io_sum = _T_43[31:0]; // @[alu.py:35:ALU.fir@42.4]
  assign io_conflag = _T_68 ? _T_46 : _T_67; // @[alu.py:44:ALU.fir@69.4]
endmodule
