module Hazard_Detection( // @[hazard_detection.py:26:Hazard_Detection.fir@2.2]
  input        clock, // @[rawmodule.py:100:Hazard_Detection.fir@3.4]
  input        reset, // @[rawmodule.py:101:Hazard_Detection.fir@4.4]
  input  [4:0] io_rs1, // @[hazard_detection.py:11:Hazard_Detection.fir@5.4]
  input  [4:0] io_rs2, // @[hazard_detection.py:11:Hazard_Detection.fir@5.4]
  input  [4:0] io_ex_rd, // @[hazard_detection.py:11:Hazard_Detection.fir@5.4]
  input  [2:0] io_Imm_Sel, // @[hazard_detection.py:11:Hazard_Detection.fir@5.4]
  input        io_ex_Mem_Read, // @[hazard_detection.py:11:Hazard_Detection.fir@5.4]
  output       io_Bubble, // @[hazard_detection.py:11:Hazard_Detection.fir@5.4]
  output       io_IF_ID_Write, // @[hazard_detection.py:11:Hazard_Detection.fir@5.4]
  output       io_PC_Write // @[hazard_detection.py:11:Hazard_Detection.fir@5.4]
);
  wire  _T_13; // @[hazard_detection.py:32:Hazard_Detection.fir@8.4]
  wire  _T_14; // @[hazard_detection.py:32:Hazard_Detection.fir@9.4]
  wire  _T_15; // @[hazard_detection.py:32:Hazard_Detection.fir@10.4]
  wire  _T_16; // @[hazard_detection.py:32:Hazard_Detection.fir@11.4]
  wire  _T_17; // @[hazard_detection.py:32:Hazard_Detection.fir@12.4]
  wire  _T_18; // @[hazard_detection.py:32:Hazard_Detection.fir@13.4]
  wire  _T_20; // @[hazard_detection.py:36:Hazard_Detection.fir@15.4]
  wire  _T_21; // @[hazard_detection.py:36:Hazard_Detection.fir@16.4]
  wire  _T_22; // @[hazard_detection.py:36:Hazard_Detection.fir@17.4]
  wire  _T_23; // @[hazard_detection.py:36:Hazard_Detection.fir@18.4]
  wire  _T_24; // @[hazard_detection.py:36:Hazard_Detection.fir@19.4]
  wire  _T_25; // @[hazard_detection.py:36:Hazard_Detection.fir@20.4]
  wire  _T_26; // @[hazard_detection.py:38:Hazard_Detection.fir@21.4]
  assign _T_13 = io_Imm_Sel == 3'h5; // @[hazard_detection.py:32:Hazard_Detection.fir@8.4]
  assign _T_14 = io_ex_Mem_Read & _T_13; // @[hazard_detection.py:32:Hazard_Detection.fir@9.4]
  assign _T_15 = io_Imm_Sel == 3'h6; // @[hazard_detection.py:32:Hazard_Detection.fir@10.4]
  assign _T_16 = _T_14 & _T_15; // @[hazard_detection.py:32:Hazard_Detection.fir@11.4]
  assign _T_17 = io_rs1 == io_ex_rd; // @[hazard_detection.py:32:Hazard_Detection.fir@12.4]
  assign _T_18 = _T_16 & _T_17; // @[hazard_detection.py:32:Hazard_Detection.fir@13.4]
  assign _T_20 = io_Imm_Sel == 3'h1; // @[hazard_detection.py:36:Hazard_Detection.fir@15.4]
  assign _T_21 = io_Imm_Sel == 3'h4; // @[hazard_detection.py:36:Hazard_Detection.fir@16.4]
  assign _T_22 = _T_20 | _T_21; // @[hazard_detection.py:36:Hazard_Detection.fir@17.4]
  assign _T_23 = io_ex_Mem_Read & _T_22; // @[hazard_detection.py:36:Hazard_Detection.fir@18.4]
  assign _T_24 = io_rs2 == io_ex_rd; // @[hazard_detection.py:36:Hazard_Detection.fir@19.4]
  assign _T_25 = _T_23 & _T_24; // @[hazard_detection.py:36:Hazard_Detection.fir@20.4]
  assign _T_26 = _T_18 | _T_25; // @[hazard_detection.py:38:Hazard_Detection.fir@21.4]
  assign io_Bubble = _T_18 | _T_25; // @[hazard_detection.py:40:Hazard_Detection.fir@23.4]
  assign io_IF_ID_Write = _T_26 ? 1'h0 : 1'h1; // @[hazard_detection.py:41:Hazard_Detection.fir@25.4]
  assign io_PC_Write = _T_26 ? 1'h0 : 1'h1; // @[hazard_detection.py:42:Hazard_Detection.fir@27.4]
endmodule
