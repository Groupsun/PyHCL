module Forward( // @[forward.py:28:Forward.fir@2.2]
  input        clock, // @[rawmodule.py:100:Forward.fir@3.4]
  input        reset, // @[rawmodule.py:101:Forward.fir@4.4]
  input        io_ex_mem_Reg_Write, // @[forward.py:11:Forward.fir@5.4]
  input  [4:0] io_ex_mem_rd, // @[forward.py:11:Forward.fir@5.4]
  input        io_ex_mem_Mem_Write, // @[forward.py:11:Forward.fir@5.4]
  input  [4:0] io_ex_mem_rs2, // @[forward.py:11:Forward.fir@5.4]
  input        io_mem_wb_Reg_Write, // @[forward.py:11:Forward.fir@5.4]
  input  [4:0] io_mem_wb_rd, // @[forward.py:11:Forward.fir@5.4]
  input  [4:0] io_id_ex_rs1, // @[forward.py:11:Forward.fir@5.4]
  input  [4:0] io_id_ex_rs2, // @[forward.py:11:Forward.fir@5.4]
  output [1:0] io_Forward_A, // @[forward.py:11:Forward.fir@5.4]
  output [1:0] io_Forward_B, // @[forward.py:11:Forward.fir@5.4]
  output       io_MemWrite_Src // @[forward.py:11:Forward.fir@5.4]
);
  wire  _T_16; // @[forward.py:31:Forward.fir@8.4]
  wire  _T_17; // @[forward.py:31:Forward.fir@9.4]
  wire  _T_18; // @[forward.py:32:Forward.fir@10.4]
  wire  _T_19; // @[forward.py:32:Forward.fir@11.4]
  wire  _T_21; // @[forward.py:34:Forward.fir@13.4]
  wire  _T_22; // @[forward.py:34:Forward.fir@14.4]
  wire  _T_23; // @[forward.py:34:Forward.fir@15.4]
  wire  _T_24; // @[forward.py:34:Forward.fir@16.4]
  wire  _T_25; // @[forward.py:34:Forward.fir@17.4]
  wire  _T_26; // @[forward.py:34:Forward.fir@18.4]
  wire  _T_30; // @[forward.py:37:Forward.fir@22.4]
  wire  _T_31; // @[forward.py:37:Forward.fir@23.4]
  wire  _T_35; // @[forward.py:39:Forward.fir@27.4]
  wire  _T_36; // @[forward.py:39:Forward.fir@28.4]
  wire  _T_37; // @[forward.py:39:Forward.fir@29.4]
  wire  _T_38; // @[forward.py:39:Forward.fir@30.4]
  wire  _T_43; // @[forward.py:45:Forward.fir@37.4]
  wire  _T_44; // @[forward.py:46:Forward.fir@38.4]
  assign _T_16 = io_ex_mem_rd != 5'h0; // @[forward.py:31:Forward.fir@8.4]
  assign _T_17 = io_ex_mem_Reg_Write & _T_16; // @[forward.py:31:Forward.fir@9.4]
  assign _T_18 = io_ex_mem_rd == io_id_ex_rs1; // @[forward.py:32:Forward.fir@10.4]
  assign _T_19 = _T_17 & _T_18; // @[forward.py:32:Forward.fir@11.4]
  assign _T_21 = io_mem_wb_rd != 5'h0; // @[forward.py:34:Forward.fir@13.4]
  assign _T_22 = io_mem_wb_Reg_Write & _T_21; // @[forward.py:34:Forward.fir@14.4]
  assign _T_23 = ~ _T_19; // @[forward.py:34:Forward.fir@15.4]
  assign _T_24 = _T_22 & _T_23; // @[forward.py:34:Forward.fir@16.4]
  assign _T_25 = io_mem_wb_rd == io_id_ex_rs1; // @[forward.py:34:Forward.fir@17.4]
  assign _T_26 = _T_24 & _T_25; // @[forward.py:34:Forward.fir@18.4]
  assign _T_30 = io_ex_mem_rd == io_id_ex_rs2; // @[forward.py:37:Forward.fir@22.4]
  assign _T_31 = _T_17 & _T_30; // @[forward.py:37:Forward.fir@23.4]
  assign _T_35 = ~ _T_31; // @[forward.py:39:Forward.fir@27.4]
  assign _T_36 = _T_22 & _T_35; // @[forward.py:39:Forward.fir@28.4]
  assign _T_37 = io_mem_wb_rd == io_id_ex_rs2; // @[forward.py:39:Forward.fir@29.4]
  assign _T_38 = _T_36 & _T_37; // @[forward.py:39:Forward.fir@30.4]
  assign _T_43 = io_mem_wb_Reg_Write & io_ex_mem_Mem_Write; // @[forward.py:45:Forward.fir@37.4]
  assign _T_44 = io_ex_mem_rs2 == io_mem_wb_rd; // @[forward.py:46:Forward.fir@38.4]
  assign io_Forward_A = {_T_19,_T_26}; // @[forward.py:41:Forward.fir@32.4]
  assign io_Forward_B = {_T_31,_T_38}; // @[forward.py:42:Forward.fir@34.4]
  assign io_MemWrite_Src = _T_43 & _T_44; // @[forward.py:48:Forward.fir@41.4]
endmodule
